module unsigned_multiplier_nl (a,
    b,
    product);
 input [7:0] a;
 input [7:0] b;
 output [15:0] product;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;

 sky130_fd_sc_hd__nand2_1 _286_ (.A(net48),
    .B(net45),
    .Y(_218_));
 sky130_fd_sc_hd__and4_1 _287_ (.A(net51),
    .B(net41),
    .C(net43),
    .D(net53),
    .X(_220_));
 sky130_fd_sc_hd__a22oi_1 _288_ (.A1(net51),
    .A2(net43),
    .B1(net53),
    .B2(net41),
    .Y(_221_));
 sky130_fd_sc_hd__and4bb_1 _289_ (.A_N(_221_),
    .B_N(_220_),
    .C(net49),
    .D(net44),
    .X(_222_));
 sky130_fd_sc_hd__or2_4 _290_ (.A(_220_),
    .B(_222_),
    .X(_223_));
 sky130_fd_sc_hd__and3_1 _291_ (.A(net48),
    .B(net45),
    .C(_223_),
    .X(_224_));
 sky130_fd_sc_hd__nand2_1 _292_ (.A(net16),
    .B(net58),
    .Y(_225_));
 sky130_fd_sc_hd__xnor2_2 _293_ (.A(_218_),
    .B(_223_),
    .Y(_226_));
 sky130_fd_sc_hd__a31o_1 _294_ (.A1(net16),
    .A2(net58),
    .A3(_226_),
    .B1(_224_),
    .X(_227_));
 sky130_fd_sc_hd__and4_1 _295_ (.A(net51),
    .B(net68),
    .C(net41),
    .D(net53),
    .X(_228_));
 sky130_fd_sc_hd__nand2_1 _296_ (.A(net49),
    .B(net43),
    .Y(_229_));
 sky130_fd_sc_hd__a22o_1 _297_ (.A1(net51),
    .A2(net41),
    .B1(net53),
    .B2(net68),
    .X(_230_));
 sky130_fd_sc_hd__and2b_1 _298_ (.A_N(_228_),
    .B(_230_),
    .X(_231_));
 sky130_fd_sc_hd__a31o_1 _299_ (.A1(net49),
    .A2(net3),
    .A3(_230_),
    .B1(_228_),
    .X(_232_));
 sky130_fd_sc_hd__and3_1 _300_ (.A(net16),
    .B(net45),
    .C(_232_),
    .X(_233_));
 sky130_fd_sc_hd__a21oi_1 _301_ (.A1(net16),
    .A2(net45),
    .B1(_232_),
    .Y(_234_));
 sky130_fd_sc_hd__nor2_1 _302_ (.A(_233_),
    .B(_234_),
    .Y(_235_));
 sky130_fd_sc_hd__a22o_1 _303_ (.A1(net51),
    .A2(net69),
    .B1(net50),
    .B2(net41),
    .X(_236_));
 sky130_fd_sc_hd__nand4_2 _304_ (.A(net51),
    .B(net69),
    .C(net50),
    .D(net42),
    .Y(_237_));
 sky130_fd_sc_hd__nand2_1 _305_ (.A(_236_),
    .B(_237_),
    .Y(_238_));
 sky130_fd_sc_hd__nand2_1 _306_ (.A(net48),
    .B(net3),
    .Y(_239_));
 sky130_fd_sc_hd__or2_1 _307_ (.A(_238_),
    .B(_239_),
    .X(_240_));
 sky130_fd_sc_hd__xor2_1 _308_ (.A(_238_),
    .B(_239_),
    .X(_241_));
 sky130_fd_sc_hd__and4_1 _309_ (.A(net34),
    .B(net36),
    .C(net33),
    .D(net56),
    .X(_242_));
 sky130_fd_sc_hd__nand2_1 _310_ (.A(net63),
    .B(net67),
    .Y(_243_));
 sky130_fd_sc_hd__a22oi_2 _311_ (.A1(net34),
    .A2(net33),
    .B1(net61),
    .B2(net36),
    .Y(_244_));
 sky130_fd_sc_hd__or3_4 _312_ (.A(_242_),
    .B(_243_),
    .C(_244_),
    .X(_245_));
 sky130_fd_sc_hd__o21bai_1 _313_ (.A1(_243_),
    .A2(_244_),
    .B1_N(_242_),
    .Y(_246_));
 sky130_fd_sc_hd__nand2_1 _314_ (.A(net54),
    .B(net67),
    .Y(_247_));
 sky130_fd_sc_hd__and4_1 _315_ (.A(net36),
    .B(net34),
    .C(net55),
    .D(net56),
    .X(_248_));
 sky130_fd_sc_hd__a22oi_2 _316_ (.A1(net63),
    .A2(net36),
    .B1(net57),
    .B2(net34),
    .Y(_249_));
 sky130_fd_sc_hd__or3_4 _317_ (.A(_248_),
    .B(_247_),
    .C(_249_),
    .X(_250_));
 sky130_fd_sc_hd__o21ai_1 _318_ (.A1(_248_),
    .A2(_249_),
    .B1(_247_),
    .Y(_251_));
 sky130_fd_sc_hd__nand3_1 _319_ (.A(_246_),
    .B(_250_),
    .C(_251_),
    .Y(_252_));
 sky130_fd_sc_hd__a21o_1 _320_ (.A1(_251_),
    .A2(_250_),
    .B1(_246_),
    .X(_253_));
 sky130_fd_sc_hd__nand3_1 _321_ (.A(_241_),
    .B(_252_),
    .C(_253_),
    .Y(_254_));
 sky130_fd_sc_hd__a21o_1 _322_ (.A1(_252_),
    .A2(_253_),
    .B1(_241_),
    .X(_255_));
 sky130_fd_sc_hd__o21ai_1 _323_ (.A1(_242_),
    .A2(_244_),
    .B1(_243_),
    .Y(_256_));
 sky130_fd_sc_hd__and4_1 _324_ (.A(net33),
    .B(net38),
    .C(net36),
    .D(net57),
    .X(_257_));
 sky130_fd_sc_hd__nand2_1 _325_ (.A(net68),
    .B(net63),
    .Y(_258_));
 sky130_fd_sc_hd__a22oi_2 _326_ (.A1(net36),
    .A2(net9),
    .B1(net57),
    .B2(net38),
    .Y(_259_));
 sky130_fd_sc_hd__or3_4 _327_ (.A(_257_),
    .B(_258_),
    .C(_259_),
    .X(_260_));
 sky130_fd_sc_hd__o21bai_1 _328_ (.A1(_258_),
    .A2(_259_),
    .B1_N(net70),
    .Y(_261_));
 sky130_fd_sc_hd__nand3_1 _329_ (.A(_245_),
    .B(_256_),
    .C(_261_),
    .Y(_262_));
 sky130_fd_sc_hd__xnor2_1 _330_ (.A(_229_),
    .B(_231_),
    .Y(_263_));
 sky130_fd_sc_hd__a21o_1 _331_ (.A1(_256_),
    .A2(_245_),
    .B1(_261_),
    .X(_264_));
 sky130_fd_sc_hd__nand3_1 _332_ (.A(_262_),
    .B(_263_),
    .C(_264_),
    .Y(_265_));
 sky130_fd_sc_hd__a21bo_1 _333_ (.A1(_263_),
    .A2(_264_),
    .B1_N(_262_),
    .X(_266_));
 sky130_fd_sc_hd__nand3_1 _334_ (.A(_254_),
    .B(_255_),
    .C(_266_),
    .Y(_267_));
 sky130_fd_sc_hd__a21o_1 _335_ (.A1(_254_),
    .A2(_255_),
    .B1(_266_),
    .X(_268_));
 sky130_fd_sc_hd__nand3_2 _336_ (.A(_235_),
    .B(_267_),
    .C(_268_),
    .Y(_269_));
 sky130_fd_sc_hd__a21o_1 _337_ (.A1(_268_),
    .A2(_267_),
    .B1(_235_),
    .X(_270_));
 sky130_fd_sc_hd__a21o_1 _338_ (.A1(_264_),
    .A2(_262_),
    .B1(_263_),
    .X(_271_));
 sky130_fd_sc_hd__o21ai_1 _339_ (.A1(net70),
    .A2(_259_),
    .B1(_258_),
    .Y(_272_));
 sky130_fd_sc_hd__and4_1 _340_ (.A(net57),
    .B(net38),
    .C(net9),
    .D(net39),
    .X(_273_));
 sky130_fd_sc_hd__nand2_2 _341_ (.A(net41),
    .B(net62),
    .Y(_274_));
 sky130_fd_sc_hd__a22oi_2 _342_ (.A1(net38),
    .A2(net9),
    .B1(net57),
    .B2(net68),
    .Y(_275_));
 sky130_fd_sc_hd__or3_4 _343_ (.A(_274_),
    .B(_273_),
    .C(_275_),
    .X(_276_));
 sky130_fd_sc_hd__o21bai_1 _344_ (.A1(_274_),
    .A2(_275_),
    .B1_N(_273_),
    .Y(_277_));
 sky130_fd_sc_hd__nand3_1 _345_ (.A(_260_),
    .B(_272_),
    .C(_277_),
    .Y(_278_));
 sky130_fd_sc_hd__o2bb2a_1 _346_ (.A1_N(net50),
    .A2_N(net44),
    .B1(_220_),
    .B2(_221_),
    .X(_279_));
 sky130_fd_sc_hd__nor2_4 _347_ (.A(_222_),
    .B(_279_),
    .Y(_280_));
 sky130_fd_sc_hd__a21o_1 _348_ (.A1(_272_),
    .A2(_260_),
    .B1(_277_),
    .X(_281_));
 sky130_fd_sc_hd__nand3_4 _349_ (.A(_278_),
    .B(_280_),
    .C(net59),
    .Y(_282_));
 sky130_fd_sc_hd__a21bo_1 _350_ (.A1(_280_),
    .A2(_281_),
    .B1_N(_278_),
    .X(_283_));
 sky130_fd_sc_hd__and3_1 _351_ (.A(_265_),
    .B(_271_),
    .C(_283_),
    .X(_284_));
 sky130_fd_sc_hd__nand3_1 _352_ (.A(_265_),
    .B(_271_),
    .C(_283_),
    .Y(_285_));
 sky130_fd_sc_hd__xnor2_2 _353_ (.A(_225_),
    .B(_226_),
    .Y(_000_));
 sky130_fd_sc_hd__a21o_1 _354_ (.A1(_271_),
    .A2(_265_),
    .B1(_283_),
    .X(_001_));
 sky130_fd_sc_hd__and3_4 _355_ (.A(_001_),
    .B(_000_),
    .C(_285_),
    .X(_002_));
 sky130_fd_sc_hd__o211ai_2 _356_ (.A1(_284_),
    .A2(_002_),
    .B1(_269_),
    .C1(_270_),
    .Y(_003_));
 sky130_fd_sc_hd__a211o_1 _357_ (.A1(_270_),
    .A2(_269_),
    .B1(_284_),
    .C1(_002_),
    .X(_004_));
 sky130_fd_sc_hd__and3_1 _358_ (.A(_227_),
    .B(_003_),
    .C(_004_),
    .X(_005_));
 sky130_fd_sc_hd__a21oi_2 _359_ (.A1(_003_),
    .A2(_004_),
    .B1(_227_),
    .Y(_006_));
 sky130_fd_sc_hd__nor2_2 _360_ (.A(_005_),
    .B(_006_),
    .Y(_007_));
 sky130_fd_sc_hd__a21oi_1 _361_ (.A1(_285_),
    .A2(_001_),
    .B1(_000_),
    .Y(_008_));
 sky130_fd_sc_hd__a21o_1 _362_ (.A1(_281_),
    .A2(_278_),
    .B1(_280_),
    .X(_009_));
 sky130_fd_sc_hd__and4_1 _363_ (.A(net39),
    .B(net41),
    .C(net33),
    .D(net56),
    .X(_010_));
 sky130_fd_sc_hd__nand2_1 _364_ (.A(net43),
    .B(net62),
    .Y(_011_));
 sky130_fd_sc_hd__a22oi_2 _365_ (.A1(net39),
    .A2(net33),
    .B1(net61),
    .B2(net41),
    .Y(_012_));
 sky130_fd_sc_hd__or3_4 _366_ (.A(_010_),
    .B(_011_),
    .C(_012_),
    .X(_013_));
 sky130_fd_sc_hd__o21bai_1 _367_ (.A1(_011_),
    .A2(_012_),
    .B1_N(_010_),
    .Y(_014_));
 sky130_fd_sc_hd__o21ai_1 _368_ (.A1(_273_),
    .A2(_275_),
    .B1(_274_),
    .Y(_015_));
 sky130_fd_sc_hd__nand3_1 _369_ (.A(_276_),
    .B(_014_),
    .C(_015_),
    .Y(_016_));
 sky130_fd_sc_hd__a21o_1 _370_ (.A1(_015_),
    .A2(_276_),
    .B1(_014_),
    .X(_017_));
 sky130_fd_sc_hd__and4_1 _371_ (.A(net52),
    .B(net3),
    .C(net45),
    .D(net54),
    .X(_018_));
 sky130_fd_sc_hd__nand4_1 _372_ (.A(net51),
    .B(net43),
    .C(net44),
    .D(net53),
    .Y(_019_));
 sky130_fd_sc_hd__a22o_1 _373_ (.A1(net51),
    .A2(net44),
    .B1(net53),
    .B2(net43),
    .X(_020_));
 sky130_fd_sc_hd__and2_1 _374_ (.A(net50),
    .B(net58),
    .X(_021_));
 sky130_fd_sc_hd__a21oi_1 _375_ (.A1(_019_),
    .A2(_020_),
    .B1(_021_),
    .Y(_022_));
 sky130_fd_sc_hd__and3_1 _376_ (.A(_019_),
    .B(_020_),
    .C(_021_),
    .X(_023_));
 sky130_fd_sc_hd__nor2_1 _377_ (.A(_022_),
    .B(_023_),
    .Y(_024_));
 sky130_fd_sc_hd__nand3_1 _378_ (.A(_016_),
    .B(_017_),
    .C(_024_),
    .Y(_025_));
 sky130_fd_sc_hd__a21bo_1 _379_ (.A1(_024_),
    .A2(_017_),
    .B1_N(_016_),
    .X(_026_));
 sky130_fd_sc_hd__nand3_4 _380_ (.A(_282_),
    .B(_009_),
    .C(_026_),
    .Y(_027_));
 sky130_fd_sc_hd__o211a_1 _381_ (.A1(_018_),
    .A2(_023_),
    .B1(net48),
    .C1(net58),
    .X(_028_));
 sky130_fd_sc_hd__a211oi_1 _382_ (.A1(net48),
    .A2(net58),
    .B1(_018_),
    .C1(_023_),
    .Y(_029_));
 sky130_fd_sc_hd__nor2_1 _383_ (.A(_028_),
    .B(_029_),
    .Y(_030_));
 sky130_fd_sc_hd__a21o_1 _384_ (.A1(_009_),
    .A2(_282_),
    .B1(_026_),
    .X(_031_));
 sky130_fd_sc_hd__nand3_4 _385_ (.A(_027_),
    .B(_030_),
    .C(_031_),
    .Y(_032_));
 sky130_fd_sc_hd__a211o_4 _386_ (.A1(_027_),
    .A2(_032_),
    .B1(_002_),
    .C1(_008_),
    .X(_033_));
 sky130_fd_sc_hd__o211ai_1 _387_ (.A1(_002_),
    .A2(_008_),
    .B1(_027_),
    .C1(_032_),
    .Y(_034_));
 sky130_fd_sc_hd__nand3_2 _388_ (.A(_028_),
    .B(_033_),
    .C(_034_),
    .Y(_035_));
 sky130_fd_sc_hd__nand2_1 _389_ (.A(_033_),
    .B(_035_),
    .Y(_036_));
 sky130_fd_sc_hd__a211o_1 _390_ (.A1(_033_),
    .A2(_035_),
    .B1(_006_),
    .C1(_005_),
    .X(_037_));
 sky130_fd_sc_hd__xnor2_2 _391_ (.A(_007_),
    .B(_036_),
    .Y(_038_));
 sky130_fd_sc_hd__o21ai_1 _392_ (.A1(_010_),
    .A2(_012_),
    .B1(_011_),
    .Y(_039_));
 sky130_fd_sc_hd__and4_1 _393_ (.A(net41),
    .B(net43),
    .C(net33),
    .D(net61),
    .X(_040_));
 sky130_fd_sc_hd__nand2_1 _394_ (.A(net44),
    .B(net11),
    .Y(_041_));
 sky130_fd_sc_hd__a22oi_1 _395_ (.A1(net41),
    .A2(net33),
    .B1(net61),
    .B2(net43),
    .Y(_042_));
 sky130_fd_sc_hd__nor2_1 _396_ (.A(_040_),
    .B(_042_),
    .Y(_043_));
 sky130_fd_sc_hd__o21bai_1 _397_ (.A1(_041_),
    .A2(_042_),
    .B1_N(_040_),
    .Y(_044_));
 sky130_fd_sc_hd__and3_1 _398_ (.A(_013_),
    .B(_039_),
    .C(_044_),
    .X(_045_));
 sky130_fd_sc_hd__a22o_1 _399_ (.A1(net44),
    .A2(net53),
    .B1(net58),
    .B2(net51),
    .X(_046_));
 sky130_fd_sc_hd__nand2_1 _400_ (.A(net53),
    .B(net1),
    .Y(_047_));
 sky130_fd_sc_hd__and4_1 _401_ (.A(net51),
    .B(net45),
    .C(net53),
    .D(net1),
    .X(_048_));
 sky130_fd_sc_hd__inv_2 _402_ (.A(_048_),
    .Y(_049_));
 sky130_fd_sc_hd__and2_1 _403_ (.A(_046_),
    .B(_049_),
    .X(_050_));
 sky130_fd_sc_hd__a21o_1 _404_ (.A1(_013_),
    .A2(_039_),
    .B1(_044_),
    .X(_051_));
 sky130_fd_sc_hd__and2b_1 _405_ (.A_N(_045_),
    .B(_051_),
    .X(_052_));
 sky130_fd_sc_hd__a21o_1 _406_ (.A1(_050_),
    .A2(_051_),
    .B1(_045_),
    .X(_053_));
 sky130_fd_sc_hd__a21o_1 _407_ (.A1(_016_),
    .A2(_017_),
    .B1(_024_),
    .X(_054_));
 sky130_fd_sc_hd__and3_4 _408_ (.A(_025_),
    .B(_053_),
    .C(_054_),
    .X(_055_));
 sky130_fd_sc_hd__a21oi_2 _409_ (.A1(_025_),
    .A2(_054_),
    .B1(_053_),
    .Y(_056_));
 sky130_fd_sc_hd__nor3_4 _410_ (.A(_049_),
    .B(_055_),
    .C(_056_),
    .Y(_057_));
 sky130_fd_sc_hd__a21o_1 _411_ (.A1(_031_),
    .A2(_027_),
    .B1(_030_),
    .X(_058_));
 sky130_fd_sc_hd__o211ai_2 _412_ (.A1(_055_),
    .A2(_057_),
    .B1(net66),
    .C1(_032_),
    .Y(_059_));
 sky130_fd_sc_hd__a21o_1 _413_ (.A1(_033_),
    .A2(_034_),
    .B1(_028_),
    .X(_060_));
 sky130_fd_sc_hd__and3b_1 _414_ (.A_N(_059_),
    .B(_060_),
    .C(_035_),
    .X(_061_));
 sky130_fd_sc_hd__a21bo_1 _415_ (.A1(_060_),
    .A2(_035_),
    .B1_N(_059_),
    .X(_062_));
 sky130_fd_sc_hd__nand2b_1 _416_ (.A_N(_061_),
    .B(_062_),
    .Y(_063_));
 sky130_fd_sc_hd__a211o_1 _417_ (.A1(_058_),
    .A2(_032_),
    .B1(_057_),
    .C1(_055_),
    .X(_064_));
 sky130_fd_sc_hd__o21a_1 _418_ (.A1(_055_),
    .A2(_056_),
    .B1(_049_),
    .X(_065_));
 sky130_fd_sc_hd__or2_4 _419_ (.A(_057_),
    .B(_065_),
    .X(_066_));
 sky130_fd_sc_hd__xor2_1 _420_ (.A(_050_),
    .B(_052_),
    .X(_067_));
 sky130_fd_sc_hd__xnor2_1 _421_ (.A(_041_),
    .B(_043_),
    .Y(_068_));
 sky130_fd_sc_hd__and4_1 _422_ (.A(net43),
    .B(net44),
    .C(net33),
    .D(net56),
    .X(_069_));
 sky130_fd_sc_hd__a22oi_1 _423_ (.A1(net43),
    .A2(net33),
    .B1(net56),
    .B2(net44),
    .Y(_070_));
 sky130_fd_sc_hd__and4bb_1 _424_ (.A_N(_069_),
    .B_N(_070_),
    .C(net55),
    .D(net58),
    .X(_071_));
 sky130_fd_sc_hd__nor2_1 _425_ (.A(_069_),
    .B(_071_),
    .Y(_072_));
 sky130_fd_sc_hd__and2b_1 _426_ (.A_N(_072_),
    .B(_068_),
    .X(_073_));
 sky130_fd_sc_hd__xnor2_1 _427_ (.A(_068_),
    .B(_072_),
    .Y(_074_));
 sky130_fd_sc_hd__and3_1 _428_ (.A(net53),
    .B(net1),
    .C(_074_),
    .X(_075_));
 sky130_fd_sc_hd__o21a_1 _429_ (.A1(_073_),
    .A2(_075_),
    .B1(_067_),
    .X(_076_));
 sky130_fd_sc_hd__inv_2 _430_ (.A(_076_),
    .Y(_077_));
 sky130_fd_sc_hd__and4b_1 _431_ (.A_N(_066_),
    .B(_064_),
    .C(_059_),
    .D(_076_),
    .X(_078_));
 sky130_fd_sc_hd__a2bb2o_4 _432_ (.A1_N(_066_),
    .A2_N(_077_),
    .B1(_059_),
    .B2(_064_),
    .X(_079_));
 sky130_fd_sc_hd__nand2b_1 _433_ (.A_N(_078_),
    .B(_079_),
    .Y(_080_));
 sky130_fd_sc_hd__nor3_1 _434_ (.A(_067_),
    .B(_073_),
    .C(_075_),
    .Y(_081_));
 sky130_fd_sc_hd__xnor2_1 _435_ (.A(_047_),
    .B(_074_),
    .Y(_082_));
 sky130_fd_sc_hd__o2bb2a_1 _436_ (.A1_N(net55),
    .A2_N(net58),
    .B1(_069_),
    .B2(_070_),
    .X(_083_));
 sky130_fd_sc_hd__nor2_1 _437_ (.A(_071_),
    .B(_083_),
    .Y(_084_));
 sky130_fd_sc_hd__and2_1 _438_ (.A(net33),
    .B(net58),
    .X(net17));
 sky130_fd_sc_hd__and3_1 _439_ (.A(net44),
    .B(net61),
    .C(net17),
    .X(_085_));
 sky130_fd_sc_hd__and2_1 _440_ (.A(_084_),
    .B(_085_),
    .X(_086_));
 sky130_fd_sc_hd__and2_1 _441_ (.A(_082_),
    .B(_086_),
    .X(_087_));
 sky130_fd_sc_hd__or3b_4 _442_ (.A(_076_),
    .B(_081_),
    .C_N(_087_),
    .X(_088_));
 sky130_fd_sc_hd__nor2_2 _443_ (.A(_066_),
    .B(_088_),
    .Y(_089_));
 sky130_fd_sc_hd__a21o_1 _444_ (.A1(_079_),
    .A2(_089_),
    .B1(_078_),
    .X(_090_));
 sky130_fd_sc_hd__a21oi_4 _445_ (.A1(_090_),
    .A2(_062_),
    .B1(_061_),
    .Y(_091_));
 sky130_fd_sc_hd__xor2_1 _446_ (.A(_038_),
    .B(net60),
    .X(net31));
 sky130_fd_sc_hd__a21bo_1 _447_ (.A1(_004_),
    .A2(_227_),
    .B1_N(_003_),
    .X(_092_));
 sky130_fd_sc_hd__nand4_2 _448_ (.A(net69),
    .B(net50),
    .C(net42),
    .D(net47),
    .Y(_093_));
 sky130_fd_sc_hd__a22o_1 _449_ (.A1(net40),
    .A2(net49),
    .B1(net42),
    .B2(net47),
    .X(_094_));
 sky130_fd_sc_hd__nand2_1 _450_ (.A(_093_),
    .B(_094_),
    .Y(_095_));
 sky130_fd_sc_hd__nand2_1 _451_ (.A(net3),
    .B(net46),
    .Y(_096_));
 sky130_fd_sc_hd__or2_1 _452_ (.A(_095_),
    .B(_096_),
    .X(_097_));
 sky130_fd_sc_hd__xor2_1 _453_ (.A(_095_),
    .B(_096_),
    .X(_098_));
 sky130_fd_sc_hd__and2_1 _454_ (.A(net52),
    .B(net38),
    .X(_099_));
 sky130_fd_sc_hd__nand4_1 _455_ (.A(net63),
    .B(net34),
    .C(net54),
    .D(net36),
    .Y(_100_));
 sky130_fd_sc_hd__a22o_1 _456_ (.A1(net63),
    .A2(net34),
    .B1(net54),
    .B2(net36),
    .X(_101_));
 sky130_fd_sc_hd__nand3_1 _457_ (.A(_099_),
    .B(_100_),
    .C(_101_),
    .Y(_102_));
 sky130_fd_sc_hd__a21o_1 _458_ (.A1(_100_),
    .A2(_101_),
    .B1(_099_),
    .X(_103_));
 sky130_fd_sc_hd__o21bai_1 _459_ (.A1(_247_),
    .A2(_249_),
    .B1_N(_248_),
    .Y(_104_));
 sky130_fd_sc_hd__nand3_1 _460_ (.A(_102_),
    .B(_103_),
    .C(_104_),
    .Y(_105_));
 sky130_fd_sc_hd__a21o_1 _461_ (.A1(_102_),
    .A2(_103_),
    .B1(_104_),
    .X(_106_));
 sky130_fd_sc_hd__nand3_1 _462_ (.A(_098_),
    .B(_105_),
    .C(_106_),
    .Y(_107_));
 sky130_fd_sc_hd__a21o_1 _463_ (.A1(_105_),
    .A2(_106_),
    .B1(_098_),
    .X(_108_));
 sky130_fd_sc_hd__a21bo_1 _464_ (.A1(_253_),
    .A2(_241_),
    .B1_N(_252_),
    .X(_109_));
 sky130_fd_sc_hd__and3_4 _465_ (.A(_107_),
    .B(_109_),
    .C(_108_),
    .X(_110_));
 sky130_fd_sc_hd__a21oi_1 _466_ (.A1(_107_),
    .A2(_108_),
    .B1(_109_),
    .Y(_111_));
 sky130_fd_sc_hd__a211oi_4 _467_ (.A1(_237_),
    .A2(_240_),
    .B1(_110_),
    .C1(_111_),
    .Y(_112_));
 sky130_fd_sc_hd__o211a_1 _468_ (.A1(_110_),
    .A2(_111_),
    .B1(_237_),
    .C1(_240_),
    .X(_113_));
 sky130_fd_sc_hd__a211o_1 _469_ (.A1(_267_),
    .A2(_269_),
    .B1(_113_),
    .C1(_112_),
    .X(_114_));
 sky130_fd_sc_hd__o211ai_1 _470_ (.A1(_112_),
    .A2(_113_),
    .B1(_267_),
    .C1(_269_),
    .Y(_115_));
 sky130_fd_sc_hd__nand3_1 _471_ (.A(_233_),
    .B(_114_),
    .C(_115_),
    .Y(_116_));
 sky130_fd_sc_hd__a21o_1 _472_ (.A1(_114_),
    .A2(_115_),
    .B1(_233_),
    .X(_117_));
 sky130_fd_sc_hd__and3_1 _473_ (.A(_092_),
    .B(_116_),
    .C(_117_),
    .X(_118_));
 sky130_fd_sc_hd__nand3_1 _474_ (.A(_092_),
    .B(_116_),
    .C(_117_),
    .Y(_119_));
 sky130_fd_sc_hd__a21oi_2 _475_ (.A1(_117_),
    .A2(_116_),
    .B1(_092_),
    .Y(_120_));
 sky130_fd_sc_hd__or2_1 _476_ (.A(_118_),
    .B(_120_),
    .X(_121_));
 sky130_fd_sc_hd__o21ai_1 _477_ (.A1(_038_),
    .A2(net60),
    .B1(_037_),
    .Y(_122_));
 sky130_fd_sc_hd__xnor2_1 _478_ (.A(_122_),
    .B(_121_),
    .Y(net32));
 sky130_fd_sc_hd__a22oi_1 _479_ (.A1(net40),
    .A2(net47),
    .B1(net46),
    .B2(net42),
    .Y(_123_));
 sky130_fd_sc_hd__nand2_1 _480_ (.A(net40),
    .B(net46),
    .Y(_124_));
 sky130_fd_sc_hd__and4_1 _481_ (.A(net40),
    .B(net42),
    .C(net47),
    .D(net46),
    .X(_125_));
 sky130_fd_sc_hd__nor2_1 _482_ (.A(_123_),
    .B(_125_),
    .Y(_126_));
 sky130_fd_sc_hd__nand4_1 _483_ (.A(net52),
    .B(net34),
    .C(net54),
    .D(net36),
    .Y(_127_));
 sky130_fd_sc_hd__a22o_1 _484_ (.A1(net34),
    .A2(net54),
    .B1(net36),
    .B2(net52),
    .X(_128_));
 sky130_fd_sc_hd__a22o_1 _485_ (.A1(net49),
    .A2(net67),
    .B1(_127_),
    .B2(_128_),
    .X(_129_));
 sky130_fd_sc_hd__nand4_1 _486_ (.A(net49),
    .B(net67),
    .C(_127_),
    .D(_128_),
    .Y(_130_));
 sky130_fd_sc_hd__a21bo_1 _487_ (.A1(_099_),
    .A2(_101_),
    .B1_N(_100_),
    .X(_131_));
 sky130_fd_sc_hd__nand3_1 _488_ (.A(_129_),
    .B(_130_),
    .C(_131_),
    .Y(_132_));
 sky130_fd_sc_hd__a21o_1 _489_ (.A1(_129_),
    .A2(_130_),
    .B1(_131_),
    .X(_133_));
 sky130_fd_sc_hd__nand3_1 _490_ (.A(_126_),
    .B(_132_),
    .C(_133_),
    .Y(_134_));
 sky130_fd_sc_hd__a21o_1 _491_ (.A1(_132_),
    .A2(_133_),
    .B1(_126_),
    .X(_135_));
 sky130_fd_sc_hd__a21bo_1 _492_ (.A1(_098_),
    .A2(_106_),
    .B1_N(_105_),
    .X(_136_));
 sky130_fd_sc_hd__and3_1 _493_ (.A(_134_),
    .B(_135_),
    .C(_136_),
    .X(_137_));
 sky130_fd_sc_hd__a21oi_1 _494_ (.A1(_134_),
    .A2(_135_),
    .B1(_136_),
    .Y(_138_));
 sky130_fd_sc_hd__a211o_1 _495_ (.A1(_093_),
    .A2(_097_),
    .B1(_137_),
    .C1(_138_),
    .X(_139_));
 sky130_fd_sc_hd__o211ai_2 _496_ (.A1(_137_),
    .A2(_138_),
    .B1(_093_),
    .C1(_097_),
    .Y(_140_));
 sky130_fd_sc_hd__o211ai_2 _497_ (.A1(_110_),
    .A2(_112_),
    .B1(_139_),
    .C1(_140_),
    .Y(_141_));
 sky130_fd_sc_hd__a211o_1 _498_ (.A1(_139_),
    .A2(_140_),
    .B1(_110_),
    .C1(_112_),
    .X(_142_));
 sky130_fd_sc_hd__nand2_1 _499_ (.A(_141_),
    .B(_142_),
    .Y(_143_));
 sky130_fd_sc_hd__and3_1 _500_ (.A(_114_),
    .B(_116_),
    .C(_143_),
    .X(_144_));
 sky130_fd_sc_hd__a21oi_1 _501_ (.A1(_114_),
    .A2(_116_),
    .B1(_143_),
    .Y(_145_));
 sky130_fd_sc_hd__nor2_1 _502_ (.A(_144_),
    .B(_145_),
    .Y(_146_));
 sky130_fd_sc_hd__nor3_4 _503_ (.A(_038_),
    .B(_091_),
    .C(_121_),
    .Y(_147_));
 sky130_fd_sc_hd__a21oi_2 _504_ (.A1(_037_),
    .A2(_119_),
    .B1(_120_),
    .Y(_148_));
 sky130_fd_sc_hd__nor2_1 _505_ (.A(_147_),
    .B(_148_),
    .Y(_149_));
 sky130_fd_sc_hd__xnor2_1 _506_ (.A(_146_),
    .B(_149_),
    .Y(net18));
 sky130_fd_sc_hd__and2b_1 _507_ (.A_N(_137_),
    .B(_139_),
    .X(_150_));
 sky130_fd_sc_hd__nand2_1 _508_ (.A(net49),
    .B(net34),
    .Y(_151_));
 sky130_fd_sc_hd__and4_1 _509_ (.A(net52),
    .B(net49),
    .C(net34),
    .D(net37),
    .X(_152_));
 sky130_fd_sc_hd__a22oi_1 _510_ (.A1(net52),
    .A2(net35),
    .B1(net37),
    .B2(net49),
    .Y(_153_));
 sky130_fd_sc_hd__o2bb2a_1 _511_ (.A1_N(net47),
    .A2_N(net67),
    .B1(_152_),
    .B2(_153_),
    .X(_154_));
 sky130_fd_sc_hd__and4bb_1 _512_ (.A_N(_152_),
    .B_N(_153_),
    .C(net47),
    .D(net6),
    .X(_155_));
 sky130_fd_sc_hd__nor2_1 _513_ (.A(_154_),
    .B(_155_),
    .Y(_156_));
 sky130_fd_sc_hd__nand2_1 _514_ (.A(_127_),
    .B(_130_),
    .Y(_157_));
 sky130_fd_sc_hd__xor2_1 _515_ (.A(_156_),
    .B(_157_),
    .X(_158_));
 sky130_fd_sc_hd__and3_1 _516_ (.A(net40),
    .B(net46),
    .C(_158_),
    .X(_159_));
 sky130_fd_sc_hd__xor2_1 _517_ (.A(_124_),
    .B(_158_),
    .X(_160_));
 sky130_fd_sc_hd__and2_1 _518_ (.A(_132_),
    .B(_134_),
    .X(_161_));
 sky130_fd_sc_hd__nor2_1 _519_ (.A(_160_),
    .B(_161_),
    .Y(_162_));
 sky130_fd_sc_hd__xor2_1 _520_ (.A(_160_),
    .B(_161_),
    .X(_163_));
 sky130_fd_sc_hd__xnor2_1 _521_ (.A(_125_),
    .B(_163_),
    .Y(_164_));
 sky130_fd_sc_hd__or2_1 _522_ (.A(_150_),
    .B(_164_),
    .X(_165_));
 sky130_fd_sc_hd__nand2_1 _523_ (.A(_150_),
    .B(_164_),
    .Y(_166_));
 sky130_fd_sc_hd__nand2_1 _524_ (.A(_165_),
    .B(_166_),
    .Y(_167_));
 sky130_fd_sc_hd__and2_1 _525_ (.A(_141_),
    .B(_167_),
    .X(_168_));
 sky130_fd_sc_hd__nor2_1 _526_ (.A(_141_),
    .B(_167_),
    .Y(_169_));
 sky130_fd_sc_hd__nor2_1 _527_ (.A(_168_),
    .B(_169_),
    .Y(_170_));
 sky130_fd_sc_hd__o21ba_1 _528_ (.A1(_144_),
    .A2(_149_),
    .B1_N(_145_),
    .X(_171_));
 sky130_fd_sc_hd__xnor2_1 _529_ (.A(_170_),
    .B(_171_),
    .Y(net19));
 sky130_fd_sc_hd__and4_1 _530_ (.A(net49),
    .B(net47),
    .C(net35),
    .D(net37),
    .X(_172_));
 sky130_fd_sc_hd__nand2_1 _531_ (.A(net47),
    .B(net37),
    .Y(_173_));
 sky130_fd_sc_hd__a21oi_1 _532_ (.A1(_151_),
    .A2(_173_),
    .B1(_172_),
    .Y(_174_));
 sky130_fd_sc_hd__nand2_1 _533_ (.A(net46),
    .B(net6),
    .Y(_175_));
 sky130_fd_sc_hd__xnor2_1 _534_ (.A(_174_),
    .B(_175_),
    .Y(_176_));
 sky130_fd_sc_hd__or2_1 _535_ (.A(_152_),
    .B(_155_),
    .X(_177_));
 sky130_fd_sc_hd__and2_1 _536_ (.A(_176_),
    .B(_177_),
    .X(_178_));
 sky130_fd_sc_hd__nor2_1 _537_ (.A(_176_),
    .B(_177_),
    .Y(_179_));
 sky130_fd_sc_hd__nor2_1 _538_ (.A(_178_),
    .B(_179_),
    .Y(_180_));
 sky130_fd_sc_hd__a21oi_1 _539_ (.A1(_156_),
    .A2(_157_),
    .B1(_159_),
    .Y(_181_));
 sky130_fd_sc_hd__xnor2_1 _540_ (.A(_180_),
    .B(_181_),
    .Y(_182_));
 sky130_fd_sc_hd__a21oi_1 _541_ (.A1(_125_),
    .A2(_163_),
    .B1(_162_),
    .Y(_183_));
 sky130_fd_sc_hd__nand2b_1 _542_ (.A_N(_183_),
    .B(_182_),
    .Y(_184_));
 sky130_fd_sc_hd__nand2b_1 _543_ (.A_N(_182_),
    .B(_183_),
    .Y(_185_));
 sky130_fd_sc_hd__nand2_1 _544_ (.A(_184_),
    .B(_185_),
    .Y(_186_));
 sky130_fd_sc_hd__nor2_1 _545_ (.A(_165_),
    .B(_186_),
    .Y(_187_));
 sky130_fd_sc_hd__or2_1 _546_ (.A(_165_),
    .B(_186_),
    .X(_188_));
 sky130_fd_sc_hd__and2_1 _547_ (.A(_165_),
    .B(_186_),
    .X(_189_));
 sky130_fd_sc_hd__nor2_1 _548_ (.A(_187_),
    .B(_189_),
    .Y(_190_));
 sky130_fd_sc_hd__a311o_1 _549_ (.A1(_145_),
    .A2(_165_),
    .A3(_166_),
    .B1(_148_),
    .C1(_169_),
    .X(_191_));
 sky130_fd_sc_hd__o21bai_1 _550_ (.A1(_144_),
    .A2(_168_),
    .B1_N(_169_),
    .Y(_192_));
 sky130_fd_sc_hd__o21ai_1 _551_ (.A1(_147_),
    .A2(_191_),
    .B1(_192_),
    .Y(_193_));
 sky130_fd_sc_hd__xnor2_1 _552_ (.A(_190_),
    .B(_193_),
    .Y(net20));
 sky130_fd_sc_hd__o21ai_1 _553_ (.A1(_189_),
    .A2(_193_),
    .B1(_188_),
    .Y(_194_));
 sky130_fd_sc_hd__a22o_1 _554_ (.A1(net47),
    .A2(net35),
    .B1(net37),
    .B2(net46),
    .X(_195_));
 sky130_fd_sc_hd__nand4_1 _555_ (.A(net47),
    .B(net46),
    .C(net35),
    .D(net37),
    .Y(_196_));
 sky130_fd_sc_hd__nand2_1 _556_ (.A(_195_),
    .B(_196_),
    .Y(_197_));
 sky130_fd_sc_hd__a31o_1 _557_ (.A1(net46),
    .A2(net6),
    .A3(_174_),
    .B1(_172_),
    .X(_198_));
 sky130_fd_sc_hd__and3_1 _558_ (.A(_195_),
    .B(_196_),
    .C(_198_),
    .X(_199_));
 sky130_fd_sc_hd__xnor2_1 _559_ (.A(_197_),
    .B(_198_),
    .Y(_200_));
 sky130_fd_sc_hd__o21bai_1 _560_ (.A1(_179_),
    .A2(_181_),
    .B1_N(_178_),
    .Y(_201_));
 sky130_fd_sc_hd__xnor2_1 _561_ (.A(_200_),
    .B(_201_),
    .Y(_202_));
 sky130_fd_sc_hd__xnor2_1 _562_ (.A(_184_),
    .B(_202_),
    .Y(_203_));
 sky130_fd_sc_hd__inv_2 _563_ (.A(_203_),
    .Y(_204_));
 sky130_fd_sc_hd__xnor2_1 _564_ (.A(_194_),
    .B(_203_),
    .Y(net21));
 sky130_fd_sc_hd__o2111a_1 _565_ (.A1(_147_),
    .A2(_191_),
    .B1(_192_),
    .C1(_204_),
    .D1(_190_),
    .X(_205_));
 sky130_fd_sc_hd__a21oi_1 _566_ (.A1(_184_),
    .A2(_188_),
    .B1(_202_),
    .Y(_206_));
 sky130_fd_sc_hd__and3_1 _567_ (.A(net46),
    .B(net35),
    .C(_173_),
    .X(_207_));
 sky130_fd_sc_hd__xor2_1 _568_ (.A(_199_),
    .B(_207_),
    .X(_208_));
 sky130_fd_sc_hd__and2_1 _569_ (.A(_200_),
    .B(_201_),
    .X(_209_));
 sky130_fd_sc_hd__xor2_1 _570_ (.A(_208_),
    .B(_209_),
    .X(_210_));
 sky130_fd_sc_hd__o21a_1 _571_ (.A1(_205_),
    .A2(_206_),
    .B1(_210_),
    .X(_211_));
 sky130_fd_sc_hd__or3_4 _572_ (.A(_206_),
    .B(_205_),
    .C(_210_),
    .X(_212_));
 sky130_fd_sc_hd__and2b_1 _573_ (.A_N(_211_),
    .B(_212_),
    .X(net22));
 sky130_fd_sc_hd__a21bo_1 _574_ (.A1(_199_),
    .A2(_207_),
    .B1_N(_196_),
    .X(_213_));
 sky130_fd_sc_hd__a211o_1 _575_ (.A1(_208_),
    .A2(_209_),
    .B1(_213_),
    .C1(_211_),
    .X(net23));
 sky130_fd_sc_hd__nand2_1 _576_ (.A(_077_),
    .B(_088_),
    .Y(_214_));
 sky130_fd_sc_hd__xnor2_1 _577_ (.A(_066_),
    .B(_214_),
    .Y(net28));
 sky130_fd_sc_hd__a22oi_1 _578_ (.A1(net44),
    .A2(net9),
    .B1(net58),
    .B2(net57),
    .Y(_215_));
 sky130_fd_sc_hd__nor2_1 _579_ (.A(_085_),
    .B(_215_),
    .Y(net24));
 sky130_fd_sc_hd__nor2_1 _580_ (.A(_084_),
    .B(_085_),
    .Y(_216_));
 sky130_fd_sc_hd__nor2_1 _581_ (.A(_086_),
    .B(_216_),
    .Y(net25));
 sky130_fd_sc_hd__nor2_1 _582_ (.A(_082_),
    .B(_086_),
    .Y(_217_));
 sky130_fd_sc_hd__nor2_1 _583_ (.A(_087_),
    .B(_217_),
    .Y(net26));
 sky130_fd_sc_hd__o21bai_1 _584_ (.A1(_076_),
    .A2(_081_),
    .B1_N(_087_),
    .Y(_219_));
 sky130_fd_sc_hd__and2_1 _585_ (.A(_088_),
    .B(_219_),
    .X(net27));
 sky130_fd_sc_hd__xnor2_1 _586_ (.A(_080_),
    .B(_089_),
    .Y(net29));
 sky130_fd_sc_hd__xnor2_1 _587_ (.A(_063_),
    .B(_090_),
    .Y(net30));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_125 ();
 sky130_fd_sc_hd__buf_1 input1 (.A(a[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(a[1]),
    .X(net2));
 sky130_fd_sc_hd__dlymetal6s2s_1 input3 (.A(a[2]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(a[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(a[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(a[5]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(a[6]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(a[7]),
    .X(net8));
 sky130_fd_sc_hd__buf_2 input9 (.A(b[0]),
    .X(net9));
 sky130_fd_sc_hd__buf_6 input10 (.A(b[1]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(b[2]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(b[3]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(b[4]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(b[5]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(b[6]),
    .X(net15));
 sky130_fd_sc_hd__dlymetal6s2s_1 input16 (.A(b[7]),
    .X(net16));
 sky130_fd_sc_hd__buf_2 output17 (.A(net17),
    .X(product[0]));
 sky130_fd_sc_hd__buf_4 output18 (.A(net18),
    .X(product[10]));
 sky130_fd_sc_hd__buf_4 output19 (.A(net19),
    .X(product[11]));
 sky130_fd_sc_hd__buf_4 output20 (.A(net20),
    .X(product[12]));
 sky130_fd_sc_hd__buf_6 output21 (.A(net21),
    .X(product[13]));
 sky130_fd_sc_hd__buf_6 output22 (.A(net22),
    .X(product[14]));
 sky130_fd_sc_hd__buf_6 output23 (.A(net23),
    .X(product[15]));
 sky130_fd_sc_hd__buf_2 output24 (.A(net24),
    .X(product[1]));
 sky130_fd_sc_hd__buf_2 output25 (.A(net25),
    .X(product[2]));
 sky130_fd_sc_hd__buf_2 output26 (.A(net26),
    .X(product[3]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(product[4]));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .X(product[5]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net29),
    .X(product[6]));
 sky130_fd_sc_hd__buf_2 output30 (.A(net30),
    .X(product[7]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .X(product[8]));
 sky130_fd_sc_hd__buf_6 output32 (.A(net32),
    .X(product[9]));
 sky130_fd_sc_hd__buf_6 fanout33 (.A(net9),
    .X(net33));
 sky130_fd_sc_hd__buf_6 fanout34 (.A(net8),
    .X(net34));
 sky130_fd_sc_hd__buf_1 fanout35 (.A(net8),
    .X(net35));
 sky130_fd_sc_hd__buf_6 fanout36 (.A(net7),
    .X(net36));
 sky130_fd_sc_hd__buf_1 fanout37 (.A(net7),
    .X(net37));
 sky130_fd_sc_hd__buf_6 fanout38 (.A(net6),
    .X(net38));
 sky130_fd_sc_hd__buf_6 fanout39 (.A(net5),
    .X(net39));
 sky130_fd_sc_hd__buf_1 fanout40 (.A(net5),
    .X(net40));
 sky130_fd_sc_hd__buf_2 fanout41 (.A(net4),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 fanout42 (.A(net4),
    .X(net42));
 sky130_fd_sc_hd__buf_4 fanout43 (.A(net3),
    .X(net43));
 sky130_fd_sc_hd__buf_2 fanout44 (.A(net45),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 fanout45 (.A(net2),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_2 fanout46 (.A(net16),
    .X(net46));
 sky130_fd_sc_hd__buf_2 fanout47 (.A(net15),
    .X(net47));
 sky130_fd_sc_hd__buf_1 fanout48 (.A(net15),
    .X(net48));
 sky130_fd_sc_hd__buf_2 fanout49 (.A(net14),
    .X(net49));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout50 (.A(net14),
    .X(net50));
 sky130_fd_sc_hd__buf_4 fanout51 (.A(net52),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 fanout52 (.A(net13),
    .X(net52));
 sky130_fd_sc_hd__buf_6 fanout53 (.A(net54),
    .X(net53));
 sky130_fd_sc_hd__buf_2 fanout54 (.A(net12),
    .X(net54));
 sky130_fd_sc_hd__buf_6 fanout55 (.A(net11),
    .X(net55));
 sky130_fd_sc_hd__buf_6 fanout56 (.A(net10),
    .X(net56));
 sky130_fd_sc_hd__buf_6 fanout57 (.A(net10),
    .X(net57));
 sky130_fd_sc_hd__buf_2 fanout58 (.A(net1),
    .X(net58));
 sky130_fd_sc_hd__buf_2 rebuffer1 (.A(_281_),
    .X(net59));
 sky130_fd_sc_hd__buf_6 rebuffer2 (.A(_091_),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 clone3 (.A(net10),
    .X(net61));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer4 (.A(net55),
    .X(net62));
 sky130_fd_sc_hd__buf_2 rebuffer5 (.A(net55),
    .X(net63));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer8 (.A(_058_),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 clone9 (.A(net6),
    .X(net67));
 sky130_fd_sc_hd__buf_6 rebuffer10 (.A(net39),
    .X(net68));
 sky130_fd_sc_hd__buf_4 rebuffer11 (.A(net68),
    .X(net69));
 sky130_fd_sc_hd__buf_1 rebuffer12 (.A(_257_),
    .X(net70));
 sky130_fd_sc_hd__fill_1 FILLER_0_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_161 ();
endmodule
