module pipelined_multiplier_nl (clk,
    reset,
    a,
    b,
    product);
 input clk;
 input reset;
 input [7:0] a;
 input [7:0] b;
 output [15:0] product;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire \a_pipe[0][0] ;
 wire \a_pipe[0][1] ;
 wire \a_pipe[0][2] ;
 wire \a_pipe[0][3] ;
 wire \a_pipe[0][4] ;
 wire \a_pipe[0][5] ;
 wire \a_pipe[0][6] ;
 wire \a_pipe[0][7] ;
 wire \b_pipe[0][0] ;
 wire \b_pipe[0][1] ;
 wire \b_pipe[0][2] ;
 wire \b_pipe[0][3] ;
 wire \b_pipe[0][4] ;
 wire \b_pipe[0][5] ;
 wire \b_pipe[0][6] ;
 wire \b_pipe[0][7] ;
 wire \partial_prod[0][0] ;
 wire \partial_prod[0][10] ;
 wire \partial_prod[0][11] ;
 wire \partial_prod[0][12] ;
 wire \partial_prod[0][13] ;
 wire \partial_prod[0][14] ;
 wire \partial_prod[0][15] ;
 wire \partial_prod[0][1] ;
 wire \partial_prod[0][2] ;
 wire \partial_prod[0][3] ;
 wire \partial_prod[0][4] ;
 wire \partial_prod[0][5] ;
 wire \partial_prod[0][6] ;
 wire \partial_prod[0][7] ;
 wire \partial_prod[0][8] ;
 wire \partial_prod[0][9] ;
 wire \partial_prod[1][0] ;
 wire \partial_prod[1][10] ;
 wire \partial_prod[1][11] ;
 wire \partial_prod[1][12] ;
 wire \partial_prod[1][13] ;
 wire \partial_prod[1][14] ;
 wire \partial_prod[1][15] ;
 wire \partial_prod[1][1] ;
 wire \partial_prod[1][2] ;
 wire \partial_prod[1][3] ;
 wire \partial_prod[1][4] ;
 wire \partial_prod[1][5] ;
 wire \partial_prod[1][6] ;
 wire \partial_prod[1][7] ;
 wire \partial_prod[1][8] ;
 wire \partial_prod[1][9] ;
 wire \partial_prod[2][0] ;
 wire \partial_prod[2][10] ;
 wire \partial_prod[2][11] ;
 wire \partial_prod[2][12] ;
 wire \partial_prod[2][13] ;
 wire \partial_prod[2][14] ;
 wire \partial_prod[2][15] ;
 wire \partial_prod[2][1] ;
 wire \partial_prod[2][2] ;
 wire \partial_prod[2][3] ;
 wire \partial_prod[2][4] ;
 wire \partial_prod[2][5] ;
 wire \partial_prod[2][6] ;
 wire \partial_prod[2][7] ;
 wire \partial_prod[2][8] ;
 wire \partial_prod[2][9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;

 sky130_fd_sc_hd__inv_2 _385_ (.A(net61),
    .Y(_016_));
 sky130_fd_sc_hd__and2_1 _386_ (.A(net45),
    .B(net58),
    .X(_000_));
 sky130_fd_sc_hd__a22oi_1 _387_ (.A1(net45),
    .A2(net56),
    .B1(net43),
    .B2(net58),
    .Y(_096_));
 sky130_fd_sc_hd__and3_1 _388_ (.A(net56),
    .B(net43),
    .C(_000_),
    .X(_097_));
 sky130_fd_sc_hd__nor2_1 _389_ (.A(_096_),
    .B(_097_),
    .Y(_001_));
 sky130_fd_sc_hd__nand2_1 _390_ (.A(net58),
    .B(\b_pipe[0][2] ),
    .Y(_098_));
 sky130_fd_sc_hd__and4_1 _391_ (.A(net45),
    .B(net56),
    .C(net43),
    .D(net54),
    .X(_099_));
 sky130_fd_sc_hd__a22o_1 _392_ (.A1(net56),
    .A2(net43),
    .B1(net54),
    .B2(net45),
    .X(_100_));
 sky130_fd_sc_hd__and2b_1 _393_ (.A_N(_099_),
    .B(_100_),
    .X(_101_));
 sky130_fd_sc_hd__xnor2_1 _394_ (.A(_098_),
    .B(_101_),
    .Y(_102_));
 sky130_fd_sc_hd__nand2_1 _395_ (.A(_097_),
    .B(_102_),
    .Y(_103_));
 sky130_fd_sc_hd__or2_1 _396_ (.A(_097_),
    .B(_102_),
    .X(_104_));
 sky130_fd_sc_hd__and2_1 _397_ (.A(_103_),
    .B(_104_),
    .X(_002_));
 sky130_fd_sc_hd__nand2_1 _398_ (.A(net56),
    .B(\b_pipe[0][2] ),
    .Y(_105_));
 sky130_fd_sc_hd__and4_1 _399_ (.A(net45),
    .B(net43),
    .C(net54),
    .D(net52),
    .X(_106_));
 sky130_fd_sc_hd__a22oi_1 _400_ (.A1(net43),
    .A2(net54),
    .B1(net52),
    .B2(net45),
    .Y(_107_));
 sky130_fd_sc_hd__nor2_1 _401_ (.A(_106_),
    .B(_107_),
    .Y(_108_));
 sky130_fd_sc_hd__xnor2_1 _402_ (.A(_105_),
    .B(_108_),
    .Y(_109_));
 sky130_fd_sc_hd__a31o_1 _403_ (.A1(net58),
    .A2(\b_pipe[0][2] ),
    .A3(_100_),
    .B1(_099_),
    .X(_110_));
 sky130_fd_sc_hd__and2_1 _404_ (.A(_109_),
    .B(_110_),
    .X(_111_));
 sky130_fd_sc_hd__xor2_1 _405_ (.A(_109_),
    .B(_110_),
    .X(_112_));
 sky130_fd_sc_hd__and3_1 _406_ (.A(net58),
    .B(net41),
    .C(_112_),
    .X(_113_));
 sky130_fd_sc_hd__a21oi_1 _407_ (.A1(net58),
    .A2(net41),
    .B1(_112_),
    .Y(_114_));
 sky130_fd_sc_hd__or2_1 _408_ (.A(_113_),
    .B(_114_),
    .X(_115_));
 sky130_fd_sc_hd__nor2_1 _409_ (.A(_103_),
    .B(_115_),
    .Y(_116_));
 sky130_fd_sc_hd__and2_1 _410_ (.A(_103_),
    .B(_115_),
    .X(_117_));
 sky130_fd_sc_hd__nor2_1 _411_ (.A(_116_),
    .B(_117_),
    .Y(_003_));
 sky130_fd_sc_hd__a22oi_1 _412_ (.A1(net56),
    .A2(net41),
    .B1(net39),
    .B2(net58),
    .Y(_118_));
 sky130_fd_sc_hd__and4_1 _413_ (.A(net58),
    .B(net56),
    .C(net41),
    .D(net39),
    .X(_119_));
 sky130_fd_sc_hd__nor2_1 _414_ (.A(_118_),
    .B(_119_),
    .Y(_120_));
 sky130_fd_sc_hd__nand2_1 _415_ (.A(net54),
    .B(\b_pipe[0][2] ),
    .Y(_121_));
 sky130_fd_sc_hd__and4_1 _416_ (.A(\b_pipe[0][0] ),
    .B(net43),
    .C(net52),
    .D(net51),
    .X(_122_));
 sky130_fd_sc_hd__a22oi_2 _417_ (.A1(net43),
    .A2(net52),
    .B1(net51),
    .B2(net45),
    .Y(_123_));
 sky130_fd_sc_hd__or3_1 _418_ (.A(_121_),
    .B(_122_),
    .C(_123_),
    .X(_124_));
 sky130_fd_sc_hd__o21ai_1 _419_ (.A1(_122_),
    .A2(_123_),
    .B1(_121_),
    .Y(_125_));
 sky130_fd_sc_hd__o21bai_1 _420_ (.A1(_105_),
    .A2(_107_),
    .B1_N(_106_),
    .Y(_126_));
 sky130_fd_sc_hd__and3_1 _421_ (.A(_124_),
    .B(_125_),
    .C(_126_),
    .X(_127_));
 sky130_fd_sc_hd__a21o_1 _422_ (.A1(_124_),
    .A2(_125_),
    .B1(_126_),
    .X(_128_));
 sky130_fd_sc_hd__nand2b_1 _423_ (.A_N(_127_),
    .B(_128_),
    .Y(_129_));
 sky130_fd_sc_hd__xnor2_1 _424_ (.A(_120_),
    .B(_129_),
    .Y(_130_));
 sky130_fd_sc_hd__o21a_1 _425_ (.A1(_111_),
    .A2(_113_),
    .B1(_130_),
    .X(_131_));
 sky130_fd_sc_hd__nor3_1 _426_ (.A(_111_),
    .B(_113_),
    .C(_130_),
    .Y(_132_));
 sky130_fd_sc_hd__nor2_1 _427_ (.A(_131_),
    .B(_132_),
    .Y(_133_));
 sky130_fd_sc_hd__and2_1 _428_ (.A(_116_),
    .B(_133_),
    .X(_134_));
 sky130_fd_sc_hd__nor2_1 _429_ (.A(_116_),
    .B(_133_),
    .Y(_135_));
 sky130_fd_sc_hd__nor2_1 _430_ (.A(_134_),
    .B(_135_),
    .Y(_004_));
 sky130_fd_sc_hd__a21o_1 _431_ (.A1(_120_),
    .A2(_128_),
    .B1(_127_),
    .X(_136_));
 sky130_fd_sc_hd__o21bai_1 _432_ (.A1(_121_),
    .A2(_123_),
    .B1_N(_122_),
    .Y(_137_));
 sky130_fd_sc_hd__nand2_1 _433_ (.A(\b_pipe[0][2] ),
    .B(net52),
    .Y(_138_));
 sky130_fd_sc_hd__and4_1 _434_ (.A(net45),
    .B(net43),
    .C(net51),
    .D(net50),
    .X(_139_));
 sky130_fd_sc_hd__a22oi_2 _435_ (.A1(net43),
    .A2(net51),
    .B1(net50),
    .B2(\b_pipe[0][0] ),
    .Y(_140_));
 sky130_fd_sc_hd__or3_1 _436_ (.A(_138_),
    .B(_139_),
    .C(_140_),
    .X(_141_));
 sky130_fd_sc_hd__o21ai_1 _437_ (.A1(_139_),
    .A2(_140_),
    .B1(_138_),
    .Y(_142_));
 sky130_fd_sc_hd__nand3_1 _438_ (.A(_137_),
    .B(_141_),
    .C(_142_),
    .Y(_143_));
 sky130_fd_sc_hd__a21o_1 _439_ (.A1(_141_),
    .A2(_142_),
    .B1(_137_),
    .X(_144_));
 sky130_fd_sc_hd__and4_1 _440_ (.A(net56),
    .B(net54),
    .C(net41),
    .D(net39),
    .X(_145_));
 sky130_fd_sc_hd__nand4_1 _441_ (.A(net56),
    .B(net54),
    .C(net41),
    .D(net39),
    .Y(_146_));
 sky130_fd_sc_hd__a22o_1 _442_ (.A1(net54),
    .A2(net41),
    .B1(net39),
    .B2(net56),
    .X(_147_));
 sky130_fd_sc_hd__and2_1 _443_ (.A(\a_pipe[0][0] ),
    .B(net38),
    .X(_148_));
 sky130_fd_sc_hd__a21oi_1 _444_ (.A1(_146_),
    .A2(_147_),
    .B1(_148_),
    .Y(_149_));
 sky130_fd_sc_hd__and3_1 _445_ (.A(_146_),
    .B(_147_),
    .C(_148_),
    .X(_150_));
 sky130_fd_sc_hd__nor2_1 _446_ (.A(_149_),
    .B(_150_),
    .Y(_151_));
 sky130_fd_sc_hd__nand3_1 _447_ (.A(_143_),
    .B(_144_),
    .C(_151_),
    .Y(_152_));
 sky130_fd_sc_hd__a21o_1 _448_ (.A1(_143_),
    .A2(_144_),
    .B1(_151_),
    .X(_153_));
 sky130_fd_sc_hd__and3_1 _449_ (.A(_136_),
    .B(_152_),
    .C(_153_),
    .X(_154_));
 sky130_fd_sc_hd__a21oi_1 _450_ (.A1(_152_),
    .A2(_153_),
    .B1(_136_),
    .Y(_155_));
 sky130_fd_sc_hd__nor3b_1 _451_ (.A(_154_),
    .B(_155_),
    .C_N(_119_),
    .Y(_156_));
 sky130_fd_sc_hd__inv_2 _452_ (.A(_156_),
    .Y(_157_));
 sky130_fd_sc_hd__o211a_1 _453_ (.A1(_145_),
    .A2(_150_),
    .B1(net58),
    .C1(net36),
    .X(_158_));
 sky130_fd_sc_hd__a211oi_1 _454_ (.A1(\a_pipe[0][0] ),
    .A2(net36),
    .B1(_145_),
    .C1(_150_),
    .Y(_159_));
 sky130_fd_sc_hd__nor2_1 _455_ (.A(_158_),
    .B(_159_),
    .Y(_160_));
 sky130_fd_sc_hd__nand2_1 _456_ (.A(net57),
    .B(net38),
    .Y(_161_));
 sky130_fd_sc_hd__and4_1 _457_ (.A(net54),
    .B(net52),
    .C(net41),
    .D(net39),
    .X(_162_));
 sky130_fd_sc_hd__a22o_1 _458_ (.A1(net52),
    .A2(net41),
    .B1(net39),
    .B2(net54),
    .X(_163_));
 sky130_fd_sc_hd__and2b_1 _459_ (.A_N(_162_),
    .B(_163_),
    .X(_164_));
 sky130_fd_sc_hd__xnor2_1 _460_ (.A(_161_),
    .B(_164_),
    .Y(_165_));
 sky130_fd_sc_hd__nand2_1 _461_ (.A(\b_pipe[0][2] ),
    .B(net51),
    .Y(_166_));
 sky130_fd_sc_hd__and2_1 _462_ (.A(net44),
    .B(net48),
    .X(_167_));
 sky130_fd_sc_hd__and4_1 _463_ (.A(\b_pipe[0][0] ),
    .B(net44),
    .C(net48),
    .D(net50),
    .X(_168_));
 sky130_fd_sc_hd__a22oi_2 _464_ (.A1(net45),
    .A2(net48),
    .B1(net50),
    .B2(net44),
    .Y(_169_));
 sky130_fd_sc_hd__or3_1 _465_ (.A(_166_),
    .B(_168_),
    .C(_169_),
    .X(_170_));
 sky130_fd_sc_hd__o21ai_1 _466_ (.A1(_168_),
    .A2(_169_),
    .B1(_166_),
    .Y(_171_));
 sky130_fd_sc_hd__o21bai_1 _467_ (.A1(_138_),
    .A2(_140_),
    .B1_N(_139_),
    .Y(_172_));
 sky130_fd_sc_hd__nand3_1 _468_ (.A(_170_),
    .B(_171_),
    .C(_172_),
    .Y(_173_));
 sky130_fd_sc_hd__a21o_1 _469_ (.A1(_170_),
    .A2(_171_),
    .B1(_172_),
    .X(_174_));
 sky130_fd_sc_hd__nand3_1 _470_ (.A(_165_),
    .B(_173_),
    .C(_174_),
    .Y(_175_));
 sky130_fd_sc_hd__a21o_1 _471_ (.A1(_173_),
    .A2(_174_),
    .B1(_165_),
    .X(_176_));
 sky130_fd_sc_hd__a21bo_1 _472_ (.A1(_144_),
    .A2(_151_),
    .B1_N(_143_),
    .X(_177_));
 sky130_fd_sc_hd__nand3_2 _473_ (.A(_175_),
    .B(_176_),
    .C(_177_),
    .Y(_178_));
 sky130_fd_sc_hd__a21o_1 _474_ (.A1(_175_),
    .A2(_176_),
    .B1(_177_),
    .X(_179_));
 sky130_fd_sc_hd__nand3_2 _475_ (.A(_160_),
    .B(_178_),
    .C(_179_),
    .Y(_180_));
 sky130_fd_sc_hd__a21o_1 _476_ (.A1(_178_),
    .A2(_179_),
    .B1(_160_),
    .X(_181_));
 sky130_fd_sc_hd__o211a_1 _477_ (.A1(_154_),
    .A2(net34),
    .B1(_180_),
    .C1(_181_),
    .X(_182_));
 sky130_fd_sc_hd__a211oi_1 _478_ (.A1(_180_),
    .A2(_181_),
    .B1(_154_),
    .C1(net34),
    .Y(_183_));
 sky130_fd_sc_hd__nor2_1 _479_ (.A(_182_),
    .B(_183_),
    .Y(_184_));
 sky130_fd_sc_hd__o21bai_1 _480_ (.A1(_154_),
    .A2(_155_),
    .B1_N(_119_),
    .Y(_185_));
 sky130_fd_sc_hd__nand3b_2 _481_ (.A_N(_156_),
    .B(_185_),
    .C(_131_),
    .Y(_186_));
 sky130_fd_sc_hd__nor3_1 _482_ (.A(_182_),
    .B(_183_),
    .C(_186_),
    .Y(_187_));
 sky130_fd_sc_hd__o21a_1 _483_ (.A1(_182_),
    .A2(_183_),
    .B1(_186_),
    .X(_188_));
 sky130_fd_sc_hd__or2_1 _484_ (.A(_187_),
    .B(_188_),
    .X(_189_));
 sky130_fd_sc_hd__a21o_1 _485_ (.A1(_157_),
    .A2(_185_),
    .B1(_131_),
    .X(_190_));
 sky130_fd_sc_hd__and3_1 _486_ (.A(_134_),
    .B(_186_),
    .C(_190_),
    .X(_191_));
 sky130_fd_sc_hd__xnor2_1 _487_ (.A(_189_),
    .B(_191_),
    .Y(_012_));
 sky130_fd_sc_hd__a31o_1 _488_ (.A1(net57),
    .A2(net38),
    .A3(_163_),
    .B1(_162_),
    .X(_192_));
 sky130_fd_sc_hd__nand2_1 _489_ (.A(net57),
    .B(net36),
    .Y(_193_));
 sky130_fd_sc_hd__xnor2_1 _490_ (.A(_192_),
    .B(_193_),
    .Y(_194_));
 sky130_fd_sc_hd__and3_1 _491_ (.A(\a_pipe[0][0] ),
    .B(net35),
    .C(_194_),
    .X(_195_));
 sky130_fd_sc_hd__a21oi_1 _492_ (.A1(net58),
    .A2(net35),
    .B1(_194_),
    .Y(_196_));
 sky130_fd_sc_hd__nor2_1 _493_ (.A(_195_),
    .B(_196_),
    .Y(_197_));
 sky130_fd_sc_hd__and4_1 _494_ (.A(net52),
    .B(net42),
    .C(net51),
    .D(net40),
    .X(_198_));
 sky130_fd_sc_hd__a22o_1 _495_ (.A1(net42),
    .A2(net51),
    .B1(net40),
    .B2(net52),
    .X(_199_));
 sky130_fd_sc_hd__and2b_1 _496_ (.A_N(_198_),
    .B(_199_),
    .X(_200_));
 sky130_fd_sc_hd__nand2_1 _497_ (.A(net55),
    .B(net38),
    .Y(_201_));
 sky130_fd_sc_hd__xnor2_1 _498_ (.A(_200_),
    .B(_201_),
    .Y(_202_));
 sky130_fd_sc_hd__and2_1 _499_ (.A(\b_pipe[0][2] ),
    .B(net50),
    .X(_203_));
 sky130_fd_sc_hd__a22o_1 _500_ (.A1(net44),
    .A2(net48),
    .B1(net46),
    .B2(net45),
    .X(_204_));
 sky130_fd_sc_hd__nand4_1 _501_ (.A(\b_pipe[0][0] ),
    .B(net44),
    .C(net48),
    .D(net46),
    .Y(_205_));
 sky130_fd_sc_hd__nand3_1 _502_ (.A(_203_),
    .B(_204_),
    .C(_205_),
    .Y(_206_));
 sky130_fd_sc_hd__a21o_1 _503_ (.A1(_204_),
    .A2(_205_),
    .B1(_203_),
    .X(_207_));
 sky130_fd_sc_hd__o21bai_1 _504_ (.A1(_166_),
    .A2(_169_),
    .B1_N(_168_),
    .Y(_208_));
 sky130_fd_sc_hd__nand3_1 _505_ (.A(_206_),
    .B(_207_),
    .C(_208_),
    .Y(_209_));
 sky130_fd_sc_hd__a21o_1 _506_ (.A1(_206_),
    .A2(_207_),
    .B1(_208_),
    .X(_210_));
 sky130_fd_sc_hd__nand3_1 _507_ (.A(_202_),
    .B(_209_),
    .C(_210_),
    .Y(_211_));
 sky130_fd_sc_hd__a21o_1 _508_ (.A1(_209_),
    .A2(_210_),
    .B1(_202_),
    .X(_212_));
 sky130_fd_sc_hd__a21bo_1 _509_ (.A1(_165_),
    .A2(_174_),
    .B1_N(_173_),
    .X(_213_));
 sky130_fd_sc_hd__nand3_1 _510_ (.A(_211_),
    .B(_212_),
    .C(_213_),
    .Y(_214_));
 sky130_fd_sc_hd__a21o_1 _511_ (.A1(_211_),
    .A2(_212_),
    .B1(_213_),
    .X(_215_));
 sky130_fd_sc_hd__and3_1 _512_ (.A(_197_),
    .B(_214_),
    .C(_215_),
    .X(_216_));
 sky130_fd_sc_hd__a21oi_1 _513_ (.A1(_214_),
    .A2(_215_),
    .B1(_197_),
    .Y(_217_));
 sky130_fd_sc_hd__a211o_1 _514_ (.A1(_178_),
    .A2(_180_),
    .B1(_216_),
    .C1(_217_),
    .X(_218_));
 sky130_fd_sc_hd__o211ai_2 _515_ (.A1(_216_),
    .A2(_217_),
    .B1(_178_),
    .C1(_180_),
    .Y(_219_));
 sky130_fd_sc_hd__nand3_1 _516_ (.A(_158_),
    .B(_218_),
    .C(_219_),
    .Y(_220_));
 sky130_fd_sc_hd__a21o_1 _517_ (.A1(_218_),
    .A2(_219_),
    .B1(_158_),
    .X(_221_));
 sky130_fd_sc_hd__a21oi_1 _518_ (.A1(_220_),
    .A2(_221_),
    .B1(_182_),
    .Y(_222_));
 sky130_fd_sc_hd__a21o_1 _519_ (.A1(_220_),
    .A2(_221_),
    .B1(_182_),
    .X(_223_));
 sky130_fd_sc_hd__and3_1 _520_ (.A(_182_),
    .B(_220_),
    .C(_221_),
    .X(_224_));
 sky130_fd_sc_hd__nor2_1 _521_ (.A(_222_),
    .B(_224_),
    .Y(_225_));
 sky130_fd_sc_hd__a41o_1 _522_ (.A1(_134_),
    .A2(_184_),
    .A3(_186_),
    .A4(_190_),
    .B1(_187_),
    .X(_226_));
 sky130_fd_sc_hd__xor2_1 _523_ (.A(_225_),
    .B(_226_),
    .X(_013_));
 sky130_fd_sc_hd__a31o_1 _524_ (.A1(net57),
    .A2(net36),
    .A3(_192_),
    .B1(_195_),
    .X(_227_));
 sky130_fd_sc_hd__a31o_1 _525_ (.A1(net55),
    .A2(net38),
    .A3(_199_),
    .B1(_198_),
    .X(_228_));
 sky130_fd_sc_hd__nand2_1 _526_ (.A(net55),
    .B(net36),
    .Y(_229_));
 sky130_fd_sc_hd__xnor2_1 _527_ (.A(_228_),
    .B(_229_),
    .Y(_230_));
 sky130_fd_sc_hd__and2_1 _528_ (.A(net57),
    .B(net35),
    .X(_231_));
 sky130_fd_sc_hd__nor2_1 _529_ (.A(_230_),
    .B(_231_),
    .Y(_232_));
 sky130_fd_sc_hd__and2_1 _530_ (.A(_230_),
    .B(_231_),
    .X(_233_));
 sky130_fd_sc_hd__or2_1 _531_ (.A(_232_),
    .B(_233_),
    .X(_234_));
 sky130_fd_sc_hd__and4_1 _532_ (.A(net41),
    .B(net51),
    .C(net39),
    .D(net50),
    .X(_235_));
 sky130_fd_sc_hd__a22o_1 _533_ (.A1(net51),
    .A2(net39),
    .B1(net50),
    .B2(net42),
    .X(_236_));
 sky130_fd_sc_hd__and2b_1 _534_ (.A_N(_235_),
    .B(_236_),
    .X(_237_));
 sky130_fd_sc_hd__nand2_1 _535_ (.A(net52),
    .B(net38),
    .Y(_238_));
 sky130_fd_sc_hd__xnor2_1 _536_ (.A(_237_),
    .B(_238_),
    .Y(_239_));
 sky130_fd_sc_hd__a22oi_1 _537_ (.A1(\b_pipe[0][2] ),
    .A2(net48),
    .B1(net46),
    .B2(net44),
    .Y(_240_));
 sky130_fd_sc_hd__nand2_1 _538_ (.A(\b_pipe[0][2] ),
    .B(net46),
    .Y(_241_));
 sky130_fd_sc_hd__a31oi_2 _539_ (.A1(\b_pipe[0][2] ),
    .A2(net46),
    .A3(_167_),
    .B1(_240_),
    .Y(_242_));
 sky130_fd_sc_hd__a21bo_1 _540_ (.A1(_203_),
    .A2(_204_),
    .B1_N(_205_),
    .X(_243_));
 sky130_fd_sc_hd__nand2_1 _541_ (.A(_242_),
    .B(_243_),
    .Y(_244_));
 sky130_fd_sc_hd__xor2_1 _542_ (.A(_242_),
    .B(_243_),
    .X(_245_));
 sky130_fd_sc_hd__xnor2_1 _543_ (.A(_239_),
    .B(_245_),
    .Y(_246_));
 sky130_fd_sc_hd__a21bo_1 _544_ (.A1(_202_),
    .A2(_210_),
    .B1_N(_209_),
    .X(_247_));
 sky130_fd_sc_hd__nand2b_1 _545_ (.A_N(_246_),
    .B(_247_),
    .Y(_248_));
 sky130_fd_sc_hd__xor2_1 _546_ (.A(_246_),
    .B(_247_),
    .X(_249_));
 sky130_fd_sc_hd__xor2_1 _547_ (.A(_234_),
    .B(_249_),
    .X(_250_));
 sky130_fd_sc_hd__a21boi_1 _548_ (.A1(_197_),
    .A2(_215_),
    .B1_N(_214_),
    .Y(_251_));
 sky130_fd_sc_hd__and2b_1 _549_ (.A_N(_251_),
    .B(_250_),
    .X(_252_));
 sky130_fd_sc_hd__xnor2_1 _550_ (.A(_250_),
    .B(_251_),
    .Y(_253_));
 sky130_fd_sc_hd__xor2_1 _551_ (.A(_227_),
    .B(_253_),
    .X(_254_));
 sky130_fd_sc_hd__a21bo_1 _552_ (.A1(_158_),
    .A2(_219_),
    .B1_N(_218_),
    .X(_255_));
 sky130_fd_sc_hd__and2_1 _553_ (.A(_254_),
    .B(_255_),
    .X(_256_));
 sky130_fd_sc_hd__or2_1 _554_ (.A(_254_),
    .B(_255_),
    .X(_257_));
 sky130_fd_sc_hd__xnor2_1 _555_ (.A(_254_),
    .B(_255_),
    .Y(_258_));
 sky130_fd_sc_hd__a21o_1 _556_ (.A1(_223_),
    .A2(_226_),
    .B1(_224_),
    .X(_259_));
 sky130_fd_sc_hd__xnor2_1 _557_ (.A(_258_),
    .B(_259_),
    .Y(_014_));
 sky130_fd_sc_hd__a21o_1 _558_ (.A1(_227_),
    .A2(_253_),
    .B1(_252_),
    .X(_260_));
 sky130_fd_sc_hd__a31o_1 _559_ (.A1(net55),
    .A2(net36),
    .A3(_228_),
    .B1(_233_),
    .X(_261_));
 sky130_fd_sc_hd__a31o_1 _560_ (.A1(net53),
    .A2(net38),
    .A3(_236_),
    .B1(_235_),
    .X(_262_));
 sky130_fd_sc_hd__nand2_1 _561_ (.A(net53),
    .B(net36),
    .Y(_263_));
 sky130_fd_sc_hd__xnor2_1 _562_ (.A(_262_),
    .B(_263_),
    .Y(_264_));
 sky130_fd_sc_hd__and2_1 _563_ (.A(net55),
    .B(net35),
    .X(_265_));
 sky130_fd_sc_hd__nor2_1 _564_ (.A(_264_),
    .B(_265_),
    .Y(_266_));
 sky130_fd_sc_hd__and2_1 _565_ (.A(_264_),
    .B(_265_),
    .X(_267_));
 sky130_fd_sc_hd__or2_1 _566_ (.A(_266_),
    .B(_267_),
    .X(_268_));
 sky130_fd_sc_hd__nor2_1 _567_ (.A(_167_),
    .B(_241_),
    .Y(_269_));
 sky130_fd_sc_hd__nand4_1 _568_ (.A(net42),
    .B(net40),
    .C(net49),
    .D(\a_pipe[0][5] ),
    .Y(_270_));
 sky130_fd_sc_hd__a22o_1 _569_ (.A1(net42),
    .A2(net49),
    .B1(\a_pipe[0][5] ),
    .B2(net39),
    .X(_271_));
 sky130_fd_sc_hd__nand2_1 _570_ (.A(_270_),
    .B(_271_),
    .Y(_272_));
 sky130_fd_sc_hd__and2_1 _571_ (.A(net51),
    .B(net38),
    .X(_273_));
 sky130_fd_sc_hd__xnor2_1 _572_ (.A(_272_),
    .B(_273_),
    .Y(_274_));
 sky130_fd_sc_hd__xnor2_1 _573_ (.A(_269_),
    .B(_274_),
    .Y(_275_));
 sky130_fd_sc_hd__a21boi_1 _574_ (.A1(_239_),
    .A2(_245_),
    .B1_N(_244_),
    .Y(_276_));
 sky130_fd_sc_hd__xnor2_1 _575_ (.A(_275_),
    .B(_276_),
    .Y(_277_));
 sky130_fd_sc_hd__xor2_1 _576_ (.A(_268_),
    .B(_277_),
    .X(_278_));
 sky130_fd_sc_hd__o21a_1 _577_ (.A1(_234_),
    .A2(_249_),
    .B1(_248_),
    .X(_279_));
 sky130_fd_sc_hd__nand2b_1 _578_ (.A_N(_279_),
    .B(_278_),
    .Y(_280_));
 sky130_fd_sc_hd__xnor2_1 _579_ (.A(_278_),
    .B(_279_),
    .Y(_281_));
 sky130_fd_sc_hd__nand2_1 _580_ (.A(_261_),
    .B(_281_),
    .Y(_282_));
 sky130_fd_sc_hd__xor2_1 _581_ (.A(_261_),
    .B(_281_),
    .X(_283_));
 sky130_fd_sc_hd__or2_1 _582_ (.A(_260_),
    .B(_283_),
    .X(_284_));
 sky130_fd_sc_hd__inv_2 _583_ (.A(_284_),
    .Y(_285_));
 sky130_fd_sc_hd__and2_1 _584_ (.A(_260_),
    .B(_283_),
    .X(_286_));
 sky130_fd_sc_hd__nor2_1 _585_ (.A(_285_),
    .B(_286_),
    .Y(_287_));
 sky130_fd_sc_hd__a21o_1 _586_ (.A1(_257_),
    .A2(_259_),
    .B1(_256_),
    .X(_288_));
 sky130_fd_sc_hd__xor2_1 _587_ (.A(_287_),
    .B(_288_),
    .X(_015_));
 sky130_fd_sc_hd__a31o_1 _588_ (.A1(net53),
    .A2(net36),
    .A3(_262_),
    .B1(_267_),
    .X(_289_));
 sky130_fd_sc_hd__a21bo_1 _589_ (.A1(_271_),
    .A2(_273_),
    .B1_N(_270_),
    .X(_290_));
 sky130_fd_sc_hd__and2_1 _590_ (.A(\a_pipe[0][4] ),
    .B(net37),
    .X(_291_));
 sky130_fd_sc_hd__nor2_1 _591_ (.A(_290_),
    .B(_291_),
    .Y(_292_));
 sky130_fd_sc_hd__and2_1 _592_ (.A(_290_),
    .B(_291_),
    .X(_293_));
 sky130_fd_sc_hd__nor2_1 _593_ (.A(_292_),
    .B(_293_),
    .Y(_294_));
 sky130_fd_sc_hd__nand2_1 _594_ (.A(net53),
    .B(net35),
    .Y(_295_));
 sky130_fd_sc_hd__xor2_1 _595_ (.A(_294_),
    .B(_295_),
    .X(_296_));
 sky130_fd_sc_hd__and4_1 _596_ (.A(net42),
    .B(net40),
    .C(net49),
    .D(net47),
    .X(_297_));
 sky130_fd_sc_hd__a22o_1 _597_ (.A1(net40),
    .A2(net49),
    .B1(net47),
    .B2(net42),
    .X(_298_));
 sky130_fd_sc_hd__nand2b_1 _598_ (.A_N(_297_),
    .B(_298_),
    .Y(_299_));
 sky130_fd_sc_hd__nand2_1 _599_ (.A(net50),
    .B(\b_pipe[0][5] ),
    .Y(_300_));
 sky130_fd_sc_hd__xor2_1 _600_ (.A(_299_),
    .B(_300_),
    .X(_301_));
 sky130_fd_sc_hd__o21bai_1 _601_ (.A1(_167_),
    .A2(_274_),
    .B1_N(_241_),
    .Y(_302_));
 sky130_fd_sc_hd__nand2b_1 _602_ (.A_N(_302_),
    .B(_301_),
    .Y(_303_));
 sky130_fd_sc_hd__and2b_1 _603_ (.A_N(_301_),
    .B(_302_),
    .X(_304_));
 sky130_fd_sc_hd__xnor2_1 _604_ (.A(_301_),
    .B(_302_),
    .Y(_305_));
 sky130_fd_sc_hd__xnor2_1 _605_ (.A(_296_),
    .B(_305_),
    .Y(_306_));
 sky130_fd_sc_hd__o32a_1 _606_ (.A1(_266_),
    .A2(_267_),
    .A3(_277_),
    .B1(_276_),
    .B2(_275_),
    .X(_307_));
 sky130_fd_sc_hd__nand2b_1 _607_ (.A_N(_307_),
    .B(_306_),
    .Y(_308_));
 sky130_fd_sc_hd__xnor2_1 _608_ (.A(_306_),
    .B(_307_),
    .Y(_309_));
 sky130_fd_sc_hd__nand2_1 _609_ (.A(_289_),
    .B(_309_),
    .Y(_310_));
 sky130_fd_sc_hd__xnor2_1 _610_ (.A(_289_),
    .B(_309_),
    .Y(_311_));
 sky130_fd_sc_hd__and3_1 _611_ (.A(_280_),
    .B(_282_),
    .C(_311_),
    .X(_312_));
 sky130_fd_sc_hd__a21oi_1 _612_ (.A1(_280_),
    .A2(_282_),
    .B1(_311_),
    .Y(_313_));
 sky130_fd_sc_hd__nor2_1 _613_ (.A(_312_),
    .B(_313_),
    .Y(_314_));
 sky130_fd_sc_hd__nor3b_1 _614_ (.A(_286_),
    .B(_258_),
    .C_N(_284_),
    .Y(_315_));
 sky130_fd_sc_hd__a21o_1 _615_ (.A1(_256_),
    .A2(_284_),
    .B1(_286_),
    .X(_316_));
 sky130_fd_sc_hd__a21oi_1 _616_ (.A1(_259_),
    .A2(_315_),
    .B1(_316_),
    .Y(_317_));
 sky130_fd_sc_hd__xnor2_1 _617_ (.A(_314_),
    .B(_317_),
    .Y(_006_));
 sky130_fd_sc_hd__a31o_1 _618_ (.A1(net53),
    .A2(\b_pipe[0][7] ),
    .A3(_294_),
    .B1(_293_),
    .X(_318_));
 sky130_fd_sc_hd__a22o_1 _619_ (.A1(net48),
    .A2(\b_pipe[0][5] ),
    .B1(net46),
    .B2(net40),
    .X(_319_));
 sky130_fd_sc_hd__and4_1 _620_ (.A(net40),
    .B(net48),
    .C(net38),
    .D(net46),
    .X(_320_));
 sky130_fd_sc_hd__inv_2 _621_ (.A(_320_),
    .Y(_321_));
 sky130_fd_sc_hd__nand2_1 _622_ (.A(_319_),
    .B(_321_),
    .Y(_322_));
 sky130_fd_sc_hd__a31o_1 _623_ (.A1(net50),
    .A2(\b_pipe[0][5] ),
    .A3(_298_),
    .B1(_297_),
    .X(_323_));
 sky130_fd_sc_hd__nand2_1 _624_ (.A(net50),
    .B(net36),
    .Y(_324_));
 sky130_fd_sc_hd__and3_1 _625_ (.A(\a_pipe[0][5] ),
    .B(net36),
    .C(_323_),
    .X(_325_));
 sky130_fd_sc_hd__xnor2_1 _626_ (.A(_323_),
    .B(_324_),
    .Y(_326_));
 sky130_fd_sc_hd__and2_1 _627_ (.A(\a_pipe[0][4] ),
    .B(\b_pipe[0][7] ),
    .X(_327_));
 sky130_fd_sc_hd__nor2_1 _628_ (.A(_326_),
    .B(_327_),
    .Y(_328_));
 sky130_fd_sc_hd__and2_1 _629_ (.A(_326_),
    .B(_327_),
    .X(_329_));
 sky130_fd_sc_hd__nor2_1 _630_ (.A(_328_),
    .B(_329_),
    .Y(_330_));
 sky130_fd_sc_hd__and3_1 _631_ (.A(_319_),
    .B(_321_),
    .C(_330_),
    .X(_331_));
 sky130_fd_sc_hd__xnor2_1 _632_ (.A(_322_),
    .B(_330_),
    .Y(_332_));
 sky130_fd_sc_hd__o21ai_1 _633_ (.A1(_296_),
    .A2(_304_),
    .B1(_303_),
    .Y(_333_));
 sky130_fd_sc_hd__nand2_1 _634_ (.A(_332_),
    .B(_333_),
    .Y(_334_));
 sky130_fd_sc_hd__xor2_1 _635_ (.A(_332_),
    .B(_333_),
    .X(_335_));
 sky130_fd_sc_hd__nand2_1 _636_ (.A(_318_),
    .B(_335_),
    .Y(_336_));
 sky130_fd_sc_hd__xnor2_1 _637_ (.A(_318_),
    .B(_335_),
    .Y(_337_));
 sky130_fd_sc_hd__a21oi_1 _638_ (.A1(_308_),
    .A2(_310_),
    .B1(_337_),
    .Y(_338_));
 sky130_fd_sc_hd__nand3_1 _639_ (.A(_308_),
    .B(_310_),
    .C(_337_),
    .Y(_339_));
 sky130_fd_sc_hd__nand2b_1 _640_ (.A_N(_338_),
    .B(_339_),
    .Y(_340_));
 sky130_fd_sc_hd__o21ba_1 _641_ (.A1(_312_),
    .A2(_317_),
    .B1_N(_313_),
    .X(_341_));
 sky130_fd_sc_hd__xor2_1 _642_ (.A(_340_),
    .B(_341_),
    .X(_007_));
 sky130_fd_sc_hd__nand2_1 _643_ (.A(\a_pipe[0][5] ),
    .B(net35),
    .Y(_342_));
 sky130_fd_sc_hd__and2_1 _644_ (.A(net48),
    .B(net37),
    .X(_343_));
 sky130_fd_sc_hd__nand2_1 _645_ (.A(net48),
    .B(net37),
    .Y(_344_));
 sky130_fd_sc_hd__mux2_1 _646_ (.A0(_344_),
    .A1(net37),
    .S(_320_),
    .X(_345_));
 sky130_fd_sc_hd__xor2_1 _647_ (.A(_342_),
    .B(_345_),
    .X(_346_));
 sky130_fd_sc_hd__and3_1 _648_ (.A(\b_pipe[0][5] ),
    .B(net47),
    .C(_346_),
    .X(_347_));
 sky130_fd_sc_hd__a21oi_1 _649_ (.A1(net38),
    .A2(net46),
    .B1(_346_),
    .Y(_348_));
 sky130_fd_sc_hd__nor2_1 _650_ (.A(_347_),
    .B(_348_),
    .Y(_349_));
 sky130_fd_sc_hd__and2_1 _651_ (.A(_331_),
    .B(_349_),
    .X(_350_));
 sky130_fd_sc_hd__xor2_1 _652_ (.A(_331_),
    .B(_349_),
    .X(_351_));
 sky130_fd_sc_hd__o21a_1 _653_ (.A1(_325_),
    .A2(_329_),
    .B1(_351_),
    .X(_352_));
 sky130_fd_sc_hd__nor3_1 _654_ (.A(_325_),
    .B(_329_),
    .C(_351_),
    .Y(_353_));
 sky130_fd_sc_hd__or2_1 _655_ (.A(_352_),
    .B(_353_),
    .X(_354_));
 sky130_fd_sc_hd__a21o_1 _656_ (.A1(_334_),
    .A2(_336_),
    .B1(_354_),
    .X(_355_));
 sky130_fd_sc_hd__inv_2 _657_ (.A(_355_),
    .Y(_356_));
 sky130_fd_sc_hd__nand3_1 _658_ (.A(_334_),
    .B(_336_),
    .C(_354_),
    .Y(_357_));
 sky130_fd_sc_hd__nand2_1 _659_ (.A(_355_),
    .B(_357_),
    .Y(_358_));
 sky130_fd_sc_hd__nand2b_1 _660_ (.A_N(_338_),
    .B(_312_),
    .Y(_359_));
 sky130_fd_sc_hd__a221o_1 _661_ (.A1(_256_),
    .A2(_284_),
    .B1(_313_),
    .B2(_339_),
    .C1(_286_),
    .X(_360_));
 sky130_fd_sc_hd__a211o_1 _662_ (.A1(_259_),
    .A2(_315_),
    .B1(_338_),
    .C1(_360_),
    .X(_361_));
 sky130_fd_sc_hd__and3_1 _663_ (.A(_339_),
    .B(_359_),
    .C(_361_),
    .X(_362_));
 sky130_fd_sc_hd__and4b_1 _664_ (.A_N(_358_),
    .B(_359_),
    .C(_361_),
    .D(_339_),
    .X(_363_));
 sky130_fd_sc_hd__xnor2_1 _665_ (.A(_358_),
    .B(_362_),
    .Y(_008_));
 sky130_fd_sc_hd__a22o_1 _666_ (.A1(net37),
    .A2(net47),
    .B1(net35),
    .B2(net49),
    .X(_364_));
 sky130_fd_sc_hd__nand3_1 _667_ (.A(net47),
    .B(net35),
    .C(_343_),
    .Y(_365_));
 sky130_fd_sc_hd__and3_1 _668_ (.A(_347_),
    .B(_364_),
    .C(_365_),
    .X(_366_));
 sky130_fd_sc_hd__a21oi_1 _669_ (.A1(_364_),
    .A2(_365_),
    .B1(_347_),
    .Y(_367_));
 sky130_fd_sc_hd__nor2_1 _670_ (.A(_366_),
    .B(_367_),
    .Y(_368_));
 sky130_fd_sc_hd__o2bb2a_1 _671_ (.A1_N(net37),
    .A2_N(_320_),
    .B1(_342_),
    .B2(_345_),
    .X(_369_));
 sky130_fd_sc_hd__and2b_1 _672_ (.A_N(_369_),
    .B(_368_),
    .X(_370_));
 sky130_fd_sc_hd__xnor2_1 _673_ (.A(_368_),
    .B(_369_),
    .Y(_371_));
 sky130_fd_sc_hd__nor3_1 _674_ (.A(_350_),
    .B(_352_),
    .C(_371_),
    .Y(_372_));
 sky130_fd_sc_hd__inv_2 _675_ (.A(_372_),
    .Y(_373_));
 sky130_fd_sc_hd__o21a_1 _676_ (.A1(_350_),
    .A2(_352_),
    .B1(_371_),
    .X(_374_));
 sky130_fd_sc_hd__o22ai_1 _677_ (.A1(_356_),
    .A2(_363_),
    .B1(_372_),
    .B2(_374_),
    .Y(_375_));
 sky130_fd_sc_hd__or4_1 _678_ (.A(_356_),
    .B(_363_),
    .C(_372_),
    .D(_374_),
    .X(_376_));
 sky130_fd_sc_hd__nand2_1 _679_ (.A(_375_),
    .B(_376_),
    .Y(_009_));
 sky130_fd_sc_hd__and3_1 _680_ (.A(net46),
    .B(net35),
    .C(_344_),
    .X(_377_));
 sky130_fd_sc_hd__nor2_1 _681_ (.A(_366_),
    .B(_370_),
    .Y(_378_));
 sky130_fd_sc_hd__xnor2_1 _682_ (.A(_377_),
    .B(_378_),
    .Y(_379_));
 sky130_fd_sc_hd__or2_1 _683_ (.A(_356_),
    .B(_374_),
    .X(_380_));
 sky130_fd_sc_hd__o21ai_1 _684_ (.A1(_363_),
    .A2(_380_),
    .B1(_373_),
    .Y(_381_));
 sky130_fd_sc_hd__o211a_1 _685_ (.A1(_363_),
    .A2(_380_),
    .B1(_379_),
    .C1(_373_),
    .X(_382_));
 sky130_fd_sc_hd__xnor2_1 _686_ (.A(_379_),
    .B(_381_),
    .Y(_010_));
 sky130_fd_sc_hd__o311a_1 _687_ (.A1(_343_),
    .A2(_366_),
    .A3(_370_),
    .B1(net35),
    .C1(net46),
    .X(_383_));
 sky130_fd_sc_hd__or2_1 _688_ (.A(_382_),
    .B(_383_),
    .X(_011_));
 sky130_fd_sc_hd__a21oi_1 _689_ (.A1(_186_),
    .A2(_190_),
    .B1(_134_),
    .Y(_384_));
 sky130_fd_sc_hd__nor2_1 _690_ (.A(_191_),
    .B(_384_),
    .Y(_005_));
 sky130_fd_sc_hd__inv_2 _691_ (.A(net62),
    .Y(_017_));
 sky130_fd_sc_hd__inv_2 _692_ (.A(net62),
    .Y(_018_));
 sky130_fd_sc_hd__inv_2 _693_ (.A(net62),
    .Y(_019_));
 sky130_fd_sc_hd__inv_2 _694_ (.A(net62),
    .Y(_020_));
 sky130_fd_sc_hd__inv_2 _695_ (.A(net63),
    .Y(_021_));
 sky130_fd_sc_hd__inv_2 _696_ (.A(net63),
    .Y(_022_));
 sky130_fd_sc_hd__inv_2 _697_ (.A(net63),
    .Y(_023_));
 sky130_fd_sc_hd__inv_2 _698_ (.A(net64),
    .Y(_024_));
 sky130_fd_sc_hd__inv_2 _699_ (.A(net64),
    .Y(_025_));
 sky130_fd_sc_hd__inv_2 _700_ (.A(net64),
    .Y(_026_));
 sky130_fd_sc_hd__inv_2 _701_ (.A(net64),
    .Y(_027_));
 sky130_fd_sc_hd__inv_2 _702_ (.A(net65),
    .Y(_028_));
 sky130_fd_sc_hd__inv_2 _703_ (.A(net65),
    .Y(_029_));
 sky130_fd_sc_hd__inv_2 _704_ (.A(net65),
    .Y(_030_));
 sky130_fd_sc_hd__inv_2 _705_ (.A(net65),
    .Y(_031_));
 sky130_fd_sc_hd__inv_2 _706_ (.A(net59),
    .Y(_032_));
 sky130_fd_sc_hd__inv_2 _707_ (.A(net59),
    .Y(_033_));
 sky130_fd_sc_hd__inv_2 _708_ (.A(net59),
    .Y(_034_));
 sky130_fd_sc_hd__inv_2 _709_ (.A(net59),
    .Y(_035_));
 sky130_fd_sc_hd__inv_2 _710_ (.A(net59),
    .Y(_036_));
 sky130_fd_sc_hd__inv_2 _711_ (.A(net60),
    .Y(_037_));
 sky130_fd_sc_hd__inv_2 _712_ (.A(net60),
    .Y(_038_));
 sky130_fd_sc_hd__inv_2 _713_ (.A(net60),
    .Y(_039_));
 sky130_fd_sc_hd__inv_2 _714_ (.A(net59),
    .Y(_040_));
 sky130_fd_sc_hd__inv_2 _715_ (.A(net59),
    .Y(_041_));
 sky130_fd_sc_hd__inv_2 _716_ (.A(net59),
    .Y(_042_));
 sky130_fd_sc_hd__inv_2 _717_ (.A(net59),
    .Y(_043_));
 sky130_fd_sc_hd__inv_2 _718_ (.A(net59),
    .Y(_044_));
 sky130_fd_sc_hd__inv_2 _719_ (.A(net60),
    .Y(_045_));
 sky130_fd_sc_hd__inv_2 _720_ (.A(net60),
    .Y(_046_));
 sky130_fd_sc_hd__inv_2 _721_ (.A(net60),
    .Y(_047_));
 sky130_fd_sc_hd__inv_2 _722_ (.A(net60),
    .Y(_048_));
 sky130_fd_sc_hd__inv_2 _723_ (.A(net60),
    .Y(_049_));
 sky130_fd_sc_hd__inv_2 _724_ (.A(net61),
    .Y(_050_));
 sky130_fd_sc_hd__inv_2 _725_ (.A(net61),
    .Y(_051_));
 sky130_fd_sc_hd__inv_2 _726_ (.A(net61),
    .Y(_052_));
 sky130_fd_sc_hd__inv_2 _727_ (.A(net61),
    .Y(_053_));
 sky130_fd_sc_hd__inv_2 _728_ (.A(net61),
    .Y(_054_));
 sky130_fd_sc_hd__inv_2 _729_ (.A(net68),
    .Y(_055_));
 sky130_fd_sc_hd__inv_2 _730_ (.A(net67),
    .Y(_056_));
 sky130_fd_sc_hd__inv_2 _731_ (.A(net67),
    .Y(_057_));
 sky130_fd_sc_hd__inv_2 _732_ (.A(net67),
    .Y(_058_));
 sky130_fd_sc_hd__inv_2 _733_ (.A(net67),
    .Y(_059_));
 sky130_fd_sc_hd__inv_2 _734_ (.A(net67),
    .Y(_060_));
 sky130_fd_sc_hd__inv_2 _735_ (.A(net67),
    .Y(_061_));
 sky130_fd_sc_hd__inv_2 _736_ (.A(net67),
    .Y(_062_));
 sky130_fd_sc_hd__inv_2 _737_ (.A(net67),
    .Y(_063_));
 sky130_fd_sc_hd__inv_2 _738_ (.A(net61),
    .Y(_064_));
 sky130_fd_sc_hd__inv_2 _739_ (.A(net61),
    .Y(_065_));
 sky130_fd_sc_hd__inv_2 _740_ (.A(net62),
    .Y(_066_));
 sky130_fd_sc_hd__inv_2 _741_ (.A(net62),
    .Y(_067_));
 sky130_fd_sc_hd__inv_2 _742_ (.A(net62),
    .Y(_068_));
 sky130_fd_sc_hd__inv_2 _743_ (.A(net63),
    .Y(_069_));
 sky130_fd_sc_hd__inv_2 _744_ (.A(net63),
    .Y(_070_));
 sky130_fd_sc_hd__inv_2 _745_ (.A(net63),
    .Y(_071_));
 sky130_fd_sc_hd__inv_2 _746_ (.A(net64),
    .Y(_072_));
 sky130_fd_sc_hd__inv_2 _747_ (.A(net64),
    .Y(_073_));
 sky130_fd_sc_hd__inv_2 _748_ (.A(net64),
    .Y(_074_));
 sky130_fd_sc_hd__inv_2 _749_ (.A(net64),
    .Y(_075_));
 sky130_fd_sc_hd__inv_2 _750_ (.A(net65),
    .Y(_076_));
 sky130_fd_sc_hd__inv_2 _751_ (.A(net65),
    .Y(_077_));
 sky130_fd_sc_hd__inv_2 _752_ (.A(net65),
    .Y(_078_));
 sky130_fd_sc_hd__inv_2 _753_ (.A(net67),
    .Y(_079_));
 sky130_fd_sc_hd__inv_2 _754_ (.A(net61),
    .Y(_080_));
 sky130_fd_sc_hd__inv_2 _755_ (.A(net61),
    .Y(_081_));
 sky130_fd_sc_hd__inv_2 _756_ (.A(net62),
    .Y(_082_));
 sky130_fd_sc_hd__inv_2 _757_ (.A(net62),
    .Y(_083_));
 sky130_fd_sc_hd__inv_2 _758_ (.A(net62),
    .Y(_084_));
 sky130_fd_sc_hd__inv_2 _759_ (.A(net63),
    .Y(_085_));
 sky130_fd_sc_hd__inv_2 _760_ (.A(net63),
    .Y(_086_));
 sky130_fd_sc_hd__inv_2 _761_ (.A(net63),
    .Y(_087_));
 sky130_fd_sc_hd__inv_2 _762_ (.A(net64),
    .Y(_088_));
 sky130_fd_sc_hd__inv_2 _763_ (.A(net64),
    .Y(_089_));
 sky130_fd_sc_hd__inv_2 _764_ (.A(net66),
    .Y(_090_));
 sky130_fd_sc_hd__inv_2 _765_ (.A(net66),
    .Y(_091_));
 sky130_fd_sc_hd__inv_2 _766_ (.A(net65),
    .Y(_092_));
 sky130_fd_sc_hd__inv_2 _767_ (.A(net65),
    .Y(_093_));
 sky130_fd_sc_hd__inv_2 _768_ (.A(net66),
    .Y(_094_));
 sky130_fd_sc_hd__inv_2 _769_ (.A(net65),
    .Y(_095_));
 sky130_fd_sc_hd__dfrtp_1 _770_ (.CLK(clknet_3_2__leaf_clk),
    .D(net92),
    .RESET_B(_016_),
    .Q(net18));
 sky130_fd_sc_hd__dfrtp_1 _771_ (.CLK(clknet_3_2__leaf_clk),
    .D(net115),
    .RESET_B(_017_),
    .Q(net25));
 sky130_fd_sc_hd__dfrtp_1 _772_ (.CLK(clknet_3_2__leaf_clk),
    .D(net110),
    .RESET_B(_018_),
    .Q(net26));
 sky130_fd_sc_hd__dfrtp_1 _773_ (.CLK(clknet_3_2__leaf_clk),
    .D(net106),
    .RESET_B(_019_),
    .Q(net27));
 sky130_fd_sc_hd__dfrtp_1 _774_ (.CLK(clknet_3_2__leaf_clk),
    .D(net89),
    .RESET_B(_020_),
    .Q(net28));
 sky130_fd_sc_hd__dfrtp_1 _775_ (.CLK(clknet_3_3__leaf_clk),
    .D(net103),
    .RESET_B(_021_),
    .Q(net29));
 sky130_fd_sc_hd__dfrtp_1 _776_ (.CLK(clknet_3_3__leaf_clk),
    .D(net102),
    .RESET_B(_022_),
    .Q(net30));
 sky130_fd_sc_hd__dfrtp_1 _777_ (.CLK(clknet_3_3__leaf_clk),
    .D(net100),
    .RESET_B(_023_),
    .Q(net31));
 sky130_fd_sc_hd__dfrtp_1 _778_ (.CLK(clknet_3_6__leaf_clk),
    .D(net85),
    .RESET_B(_024_),
    .Q(net32));
 sky130_fd_sc_hd__dfrtp_1 _779_ (.CLK(clknet_3_6__leaf_clk),
    .D(net94),
    .RESET_B(_025_),
    .Q(net33));
 sky130_fd_sc_hd__dfrtp_1 _780_ (.CLK(clknet_3_6__leaf_clk),
    .D(net108),
    .RESET_B(_026_),
    .Q(net19));
 sky130_fd_sc_hd__dfrtp_1 _781_ (.CLK(clknet_3_7__leaf_clk),
    .D(net90),
    .RESET_B(_027_),
    .Q(net20));
 sky130_fd_sc_hd__dfrtp_1 _782_ (.CLK(clknet_3_7__leaf_clk),
    .D(net97),
    .RESET_B(_028_),
    .Q(net21));
 sky130_fd_sc_hd__dfrtp_1 _783_ (.CLK(clknet_3_7__leaf_clk),
    .D(net101),
    .RESET_B(_029_),
    .Q(net22));
 sky130_fd_sc_hd__dfrtp_1 _784_ (.CLK(clknet_3_7__leaf_clk),
    .D(net98),
    .RESET_B(_030_),
    .Q(net23));
 sky130_fd_sc_hd__dfrtp_1 _785_ (.CLK(clknet_3_7__leaf_clk),
    .D(net88),
    .RESET_B(_031_),
    .Q(net24));
 sky130_fd_sc_hd__dfrtp_1 _786_ (.CLK(clknet_3_1__leaf_clk),
    .D(net1),
    .RESET_B(_032_),
    .Q(\a_pipe[0][0] ));
 sky130_fd_sc_hd__dfrtp_1 _787_ (.CLK(clknet_3_1__leaf_clk),
    .D(net2),
    .RESET_B(_033_),
    .Q(\a_pipe[0][1] ));
 sky130_fd_sc_hd__dfrtp_1 _788_ (.CLK(clknet_3_1__leaf_clk),
    .D(net3),
    .RESET_B(_034_),
    .Q(\a_pipe[0][2] ));
 sky130_fd_sc_hd__dfrtp_1 _789_ (.CLK(clknet_3_1__leaf_clk),
    .D(net4),
    .RESET_B(_035_),
    .Q(\a_pipe[0][3] ));
 sky130_fd_sc_hd__dfrtp_1 _790_ (.CLK(clknet_3_1__leaf_clk),
    .D(net5),
    .RESET_B(_036_),
    .Q(\a_pipe[0][4] ));
 sky130_fd_sc_hd__dfrtp_1 _791_ (.CLK(clknet_3_5__leaf_clk),
    .D(net6),
    .RESET_B(_037_),
    .Q(\a_pipe[0][5] ));
 sky130_fd_sc_hd__dfrtp_1 _792_ (.CLK(clknet_3_5__leaf_clk),
    .D(net7),
    .RESET_B(_038_),
    .Q(\a_pipe[0][6] ));
 sky130_fd_sc_hd__dfrtp_1 _793_ (.CLK(clknet_3_5__leaf_clk),
    .D(net8),
    .RESET_B(_039_),
    .Q(\a_pipe[0][7] ));
 sky130_fd_sc_hd__dfrtp_1 _794_ (.CLK(clknet_3_1__leaf_clk),
    .D(net9),
    .RESET_B(_040_),
    .Q(\b_pipe[0][0] ));
 sky130_fd_sc_hd__dfrtp_1 _795_ (.CLK(clknet_3_1__leaf_clk),
    .D(net10),
    .RESET_B(_041_),
    .Q(\b_pipe[0][1] ));
 sky130_fd_sc_hd__dfrtp_4 _796_ (.CLK(clknet_3_1__leaf_clk),
    .D(net11),
    .RESET_B(_042_),
    .Q(\b_pipe[0][2] ));
 sky130_fd_sc_hd__dfrtp_1 _797_ (.CLK(clknet_3_1__leaf_clk),
    .D(net12),
    .RESET_B(_043_),
    .Q(\b_pipe[0][3] ));
 sky130_fd_sc_hd__dfrtp_1 _798_ (.CLK(clknet_3_1__leaf_clk),
    .D(net13),
    .RESET_B(_044_),
    .Q(\b_pipe[0][4] ));
 sky130_fd_sc_hd__dfrtp_1 _799_ (.CLK(clknet_3_5__leaf_clk),
    .D(net14),
    .RESET_B(_045_),
    .Q(\b_pipe[0][5] ));
 sky130_fd_sc_hd__dfrtp_1 _800_ (.CLK(clknet_3_5__leaf_clk),
    .D(net15),
    .RESET_B(_046_),
    .Q(\b_pipe[0][6] ));
 sky130_fd_sc_hd__dfrtp_1 _801_ (.CLK(clknet_3_5__leaf_clk),
    .D(net16),
    .RESET_B(_047_),
    .Q(\b_pipe[0][7] ));
 sky130_fd_sc_hd__dfrtp_1 _802_ (.CLK(clknet_3_0__leaf_clk),
    .D(_000_),
    .RESET_B(_048_),
    .Q(\partial_prod[0][0] ));
 sky130_fd_sc_hd__dfrtp_1 _803_ (.CLK(clknet_3_0__leaf_clk),
    .D(_001_),
    .RESET_B(_049_),
    .Q(\partial_prod[0][1] ));
 sky130_fd_sc_hd__dfrtp_1 _804_ (.CLK(clknet_3_2__leaf_clk),
    .D(_002_),
    .RESET_B(_050_),
    .Q(\partial_prod[0][2] ));
 sky130_fd_sc_hd__dfrtp_1 _805_ (.CLK(clknet_3_0__leaf_clk),
    .D(_003_),
    .RESET_B(_051_),
    .Q(\partial_prod[0][3] ));
 sky130_fd_sc_hd__dfrtp_1 _806_ (.CLK(clknet_3_0__leaf_clk),
    .D(_004_),
    .RESET_B(_052_),
    .Q(\partial_prod[0][4] ));
 sky130_fd_sc_hd__dfrtp_1 _807_ (.CLK(clknet_3_0__leaf_clk),
    .D(_005_),
    .RESET_B(_053_),
    .Q(\partial_prod[0][5] ));
 sky130_fd_sc_hd__dfrtp_1 _808_ (.CLK(clknet_3_3__leaf_clk),
    .D(_012_),
    .RESET_B(_054_),
    .Q(\partial_prod[0][6] ));
 sky130_fd_sc_hd__dfrtp_1 _809_ (.CLK(clknet_3_3__leaf_clk),
    .D(_013_),
    .RESET_B(_055_),
    .Q(\partial_prod[0][7] ));
 sky130_fd_sc_hd__dfrtp_1 _810_ (.CLK(clknet_3_6__leaf_clk),
    .D(_014_),
    .RESET_B(_056_),
    .Q(\partial_prod[0][8] ));
 sky130_fd_sc_hd__dfrtp_1 _811_ (.CLK(clknet_3_4__leaf_clk),
    .D(_015_),
    .RESET_B(_057_),
    .Q(\partial_prod[0][9] ));
 sky130_fd_sc_hd__dfrtp_1 _812_ (.CLK(clknet_3_4__leaf_clk),
    .D(_006_),
    .RESET_B(_058_),
    .Q(\partial_prod[0][10] ));
 sky130_fd_sc_hd__dfrtp_1 _813_ (.CLK(clknet_3_4__leaf_clk),
    .D(_007_),
    .RESET_B(_059_),
    .Q(\partial_prod[0][11] ));
 sky130_fd_sc_hd__dfrtp_1 _814_ (.CLK(clknet_3_4__leaf_clk),
    .D(_008_),
    .RESET_B(_060_),
    .Q(\partial_prod[0][12] ));
 sky130_fd_sc_hd__dfrtp_1 _815_ (.CLK(clknet_3_5__leaf_clk),
    .D(_009_),
    .RESET_B(_061_),
    .Q(\partial_prod[0][13] ));
 sky130_fd_sc_hd__dfrtp_1 _816_ (.CLK(clknet_3_4__leaf_clk),
    .D(_010_),
    .RESET_B(_062_),
    .Q(\partial_prod[0][14] ));
 sky130_fd_sc_hd__dfrtp_1 _817_ (.CLK(clknet_3_4__leaf_clk),
    .D(_011_),
    .RESET_B(_063_),
    .Q(\partial_prod[0][15] ));
 sky130_fd_sc_hd__dfrtp_1 _818_ (.CLK(clknet_3_0__leaf_clk),
    .D(net111),
    .RESET_B(_064_),
    .Q(\partial_prod[1][0] ));
 sky130_fd_sc_hd__dfrtp_1 _819_ (.CLK(clknet_3_0__leaf_clk),
    .D(net80),
    .RESET_B(_065_),
    .Q(\partial_prod[1][1] ));
 sky130_fd_sc_hd__dfrtp_1 _820_ (.CLK(clknet_3_2__leaf_clk),
    .D(net114),
    .RESET_B(_066_),
    .Q(\partial_prod[1][2] ));
 sky130_fd_sc_hd__dfrtp_1 _821_ (.CLK(clknet_3_3__leaf_clk),
    .D(net83),
    .RESET_B(_067_),
    .Q(\partial_prod[1][3] ));
 sky130_fd_sc_hd__dfrtp_1 _822_ (.CLK(clknet_3_3__leaf_clk),
    .D(net75),
    .RESET_B(_068_),
    .Q(\partial_prod[1][4] ));
 sky130_fd_sc_hd__dfrtp_1 _823_ (.CLK(clknet_3_3__leaf_clk),
    .D(net77),
    .RESET_B(_069_),
    .Q(\partial_prod[1][5] ));
 sky130_fd_sc_hd__dfrtp_1 _824_ (.CLK(clknet_3_3__leaf_clk),
    .D(net109),
    .RESET_B(_070_),
    .Q(\partial_prod[1][6] ));
 sky130_fd_sc_hd__dfrtp_1 _825_ (.CLK(clknet_3_3__leaf_clk),
    .D(net104),
    .RESET_B(_071_),
    .Q(\partial_prod[1][7] ));
 sky130_fd_sc_hd__dfrtp_1 _826_ (.CLK(clknet_3_6__leaf_clk),
    .D(net79),
    .RESET_B(_072_),
    .Q(\partial_prod[1][8] ));
 sky130_fd_sc_hd__dfrtp_1 _827_ (.CLK(clknet_3_6__leaf_clk),
    .D(net84),
    .RESET_B(_073_),
    .Q(\partial_prod[1][9] ));
 sky130_fd_sc_hd__dfrtp_1 _828_ (.CLK(clknet_3_7__leaf_clk),
    .D(net73),
    .RESET_B(_074_),
    .Q(\partial_prod[1][10] ));
 sky130_fd_sc_hd__dfrtp_1 _829_ (.CLK(clknet_3_4__leaf_clk),
    .D(net95),
    .RESET_B(_075_),
    .Q(\partial_prod[1][11] ));
 sky130_fd_sc_hd__dfrtp_1 _830_ (.CLK(clknet_3_4__leaf_clk),
    .D(net82),
    .RESET_B(_076_),
    .Q(\partial_prod[1][12] ));
 sky130_fd_sc_hd__dfrtp_1 _831_ (.CLK(clknet_3_7__leaf_clk),
    .D(net113),
    .RESET_B(_077_),
    .Q(\partial_prod[1][13] ));
 sky130_fd_sc_hd__dfrtp_1 _832_ (.CLK(clknet_3_7__leaf_clk),
    .D(net71),
    .RESET_B(_078_),
    .Q(\partial_prod[1][14] ));
 sky130_fd_sc_hd__dfrtp_1 _833_ (.CLK(clknet_3_4__leaf_clk),
    .D(net91),
    .RESET_B(_079_),
    .Q(\partial_prod[1][15] ));
 sky130_fd_sc_hd__dfrtp_1 _834_ (.CLK(clknet_3_2__leaf_clk),
    .D(net70),
    .RESET_B(_080_),
    .Q(\partial_prod[2][0] ));
 sky130_fd_sc_hd__dfrtp_1 _835_ (.CLK(clknet_3_2__leaf_clk),
    .D(net69),
    .RESET_B(_081_),
    .Q(\partial_prod[2][1] ));
 sky130_fd_sc_hd__dfrtp_1 _836_ (.CLK(clknet_3_2__leaf_clk),
    .D(net112),
    .RESET_B(_082_),
    .Q(\partial_prod[2][2] ));
 sky130_fd_sc_hd__dfrtp_1 _837_ (.CLK(clknet_3_2__leaf_clk),
    .D(net81),
    .RESET_B(_083_),
    .Q(\partial_prod[2][3] ));
 sky130_fd_sc_hd__dfrtp_1 _838_ (.CLK(clknet_3_2__leaf_clk),
    .D(net107),
    .RESET_B(_084_),
    .Q(\partial_prod[2][4] ));
 sky130_fd_sc_hd__dfrtp_1 _839_ (.CLK(clknet_3_3__leaf_clk),
    .D(net87),
    .RESET_B(_085_),
    .Q(\partial_prod[2][5] ));
 sky130_fd_sc_hd__dfrtp_1 _840_ (.CLK(clknet_3_3__leaf_clk),
    .D(net99),
    .RESET_B(_086_),
    .Q(\partial_prod[2][6] ));
 sky130_fd_sc_hd__dfrtp_1 _841_ (.CLK(clknet_3_3__leaf_clk),
    .D(net86),
    .RESET_B(_087_),
    .Q(\partial_prod[2][7] ));
 sky130_fd_sc_hd__dfrtp_1 _842_ (.CLK(clknet_3_6__leaf_clk),
    .D(net96),
    .RESET_B(_088_),
    .Q(\partial_prod[2][8] ));
 sky130_fd_sc_hd__dfrtp_1 _843_ (.CLK(clknet_3_6__leaf_clk),
    .D(net78),
    .RESET_B(_089_),
    .Q(\partial_prod[2][9] ));
 sky130_fd_sc_hd__dfrtp_1 _844_ (.CLK(clknet_3_6__leaf_clk),
    .D(net116),
    .RESET_B(_090_),
    .Q(\partial_prod[2][10] ));
 sky130_fd_sc_hd__dfrtp_1 _845_ (.CLK(clknet_3_7__leaf_clk),
    .D(net76),
    .RESET_B(_091_),
    .Q(\partial_prod[2][11] ));
 sky130_fd_sc_hd__dfrtp_1 _846_ (.CLK(clknet_3_7__leaf_clk),
    .D(net74),
    .RESET_B(_092_),
    .Q(\partial_prod[2][12] ));
 sky130_fd_sc_hd__dfrtp_1 _847_ (.CLK(clknet_3_7__leaf_clk),
    .D(net93),
    .RESET_B(_093_),
    .Q(\partial_prod[2][13] ));
 sky130_fd_sc_hd__dfrtp_1 _848_ (.CLK(clknet_3_7__leaf_clk),
    .D(net105),
    .RESET_B(_094_),
    .Q(\partial_prod[2][14] ));
 sky130_fd_sc_hd__dfrtp_1 _849_ (.CLK(clknet_3_7__leaf_clk),
    .D(net72),
    .RESET_B(_095_),
    .Q(\partial_prod[2][15] ));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_215 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(a[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(a[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(a[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(a[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(a[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(a[5]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(a[6]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(a[7]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(b[0]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(b[1]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(b[2]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(b[3]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(b[4]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(b[5]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(b[6]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(b[7]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input17 (.A(reset),
    .X(net17));
 sky130_fd_sc_hd__buf_2 output18 (.A(net18),
    .X(product[0]));
 sky130_fd_sc_hd__buf_2 output19 (.A(net19),
    .X(product[10]));
 sky130_fd_sc_hd__buf_2 output20 (.A(net20),
    .X(product[11]));
 sky130_fd_sc_hd__buf_2 output21 (.A(net21),
    .X(product[12]));
 sky130_fd_sc_hd__buf_2 output22 (.A(net22),
    .X(product[13]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .X(product[14]));
 sky130_fd_sc_hd__buf_2 output24 (.A(net24),
    .X(product[15]));
 sky130_fd_sc_hd__buf_2 output25 (.A(net25),
    .X(product[1]));
 sky130_fd_sc_hd__buf_2 output26 (.A(net26),
    .X(product[2]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(product[3]));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .X(product[4]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net29),
    .X(product[5]));
 sky130_fd_sc_hd__buf_2 output30 (.A(net30),
    .X(product[6]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .X(product[7]));
 sky130_fd_sc_hd__buf_2 output32 (.A(net32),
    .X(product[8]));
 sky130_fd_sc_hd__buf_2 output33 (.A(net33),
    .X(product[9]));
 sky130_fd_sc_hd__clkbuf_1 max_cap34 (.A(_156_),
    .X(net34));
 sky130_fd_sc_hd__buf_2 fanout35 (.A(\b_pipe[0][7] ),
    .X(net35));
 sky130_fd_sc_hd__buf_2 fanout36 (.A(\b_pipe[0][6] ),
    .X(net36));
 sky130_fd_sc_hd__buf_1 fanout37 (.A(\b_pipe[0][6] ),
    .X(net37));
 sky130_fd_sc_hd__buf_2 fanout38 (.A(\b_pipe[0][5] ),
    .X(net38));
 sky130_fd_sc_hd__buf_2 fanout39 (.A(\b_pipe[0][4] ),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 fanout40 (.A(\b_pipe[0][4] ),
    .X(net40));
 sky130_fd_sc_hd__buf_2 fanout41 (.A(\b_pipe[0][3] ),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 fanout42 (.A(\b_pipe[0][3] ),
    .X(net42));
 sky130_fd_sc_hd__buf_2 fanout43 (.A(\b_pipe[0][1] ),
    .X(net43));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout44 (.A(\b_pipe[0][1] ),
    .X(net44));
 sky130_fd_sc_hd__buf_2 fanout45 (.A(\b_pipe[0][0] ),
    .X(net45));
 sky130_fd_sc_hd__buf_2 fanout46 (.A(\a_pipe[0][7] ),
    .X(net46));
 sky130_fd_sc_hd__buf_1 fanout47 (.A(\a_pipe[0][7] ),
    .X(net47));
 sky130_fd_sc_hd__buf_2 fanout48 (.A(\a_pipe[0][6] ),
    .X(net48));
 sky130_fd_sc_hd__buf_1 fanout49 (.A(\a_pipe[0][6] ),
    .X(net49));
 sky130_fd_sc_hd__buf_2 fanout50 (.A(\a_pipe[0][5] ),
    .X(net50));
 sky130_fd_sc_hd__buf_2 fanout51 (.A(\a_pipe[0][4] ),
    .X(net51));
 sky130_fd_sc_hd__buf_2 fanout52 (.A(\a_pipe[0][3] ),
    .X(net52));
 sky130_fd_sc_hd__buf_1 fanout53 (.A(\a_pipe[0][3] ),
    .X(net53));
 sky130_fd_sc_hd__buf_2 fanout54 (.A(\a_pipe[0][2] ),
    .X(net54));
 sky130_fd_sc_hd__buf_1 fanout55 (.A(\a_pipe[0][2] ),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 fanout56 (.A(\a_pipe[0][1] ),
    .X(net56));
 sky130_fd_sc_hd__buf_1 fanout57 (.A(\a_pipe[0][1] ),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 fanout58 (.A(\a_pipe[0][0] ),
    .X(net58));
 sky130_fd_sc_hd__buf_4 fanout59 (.A(net60),
    .X(net59));
 sky130_fd_sc_hd__buf_4 fanout60 (.A(net17),
    .X(net60));
 sky130_fd_sc_hd__buf_4 fanout61 (.A(net68),
    .X(net61));
 sky130_fd_sc_hd__buf_4 fanout62 (.A(net68),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_4 fanout63 (.A(net68),
    .X(net63));
 sky130_fd_sc_hd__buf_4 fanout64 (.A(net66),
    .X(net64));
 sky130_fd_sc_hd__buf_4 fanout65 (.A(net66),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_2 fanout66 (.A(net67),
    .X(net66));
 sky130_fd_sc_hd__buf_4 fanout67 (.A(net68),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_2 fanout68 (.A(net17),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__clkinv_4 clkload0 (.A(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkinv_2 clkload1 (.A(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload2 (.A(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__bufinv_16 clkload3 (.A(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkinv_4 clkload4 (.A(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__bufinv_16 clkload5 (.A(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\partial_prod[1][1] ),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\partial_prod[1][0] ),
    .X(net70));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\partial_prod[0][14] ),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\partial_prod[1][15] ),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\partial_prod[0][10] ),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\partial_prod[1][12] ),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\partial_prod[0][4] ),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\partial_prod[1][11] ),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\partial_prod[0][5] ),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\partial_prod[1][9] ),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\partial_prod[0][8] ),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\partial_prod[0][1] ),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\partial_prod[1][3] ),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\partial_prod[0][12] ),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\partial_prod[0][3] ),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\partial_prod[0][9] ),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\partial_prod[2][8] ),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\partial_prod[1][7] ),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\partial_prod[1][5] ),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\partial_prod[2][15] ),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\partial_prod[2][4] ),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\partial_prod[2][11] ),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\partial_prod[0][15] ),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\partial_prod[2][0] ),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\partial_prod[1][13] ),
    .X(net93));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\partial_prod[2][9] ),
    .X(net94));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\partial_prod[0][11] ),
    .X(net95));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\partial_prod[1][8] ),
    .X(net96));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\partial_prod[2][12] ),
    .X(net97));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\partial_prod[2][14] ),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\partial_prod[1][6] ),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\partial_prod[2][7] ),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\partial_prod[2][13] ),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\partial_prod[2][6] ),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\partial_prod[2][5] ),
    .X(net103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\partial_prod[0][7] ),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\partial_prod[1][14] ),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\partial_prod[2][3] ),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\partial_prod[1][4] ),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\partial_prod[2][10] ),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\partial_prod[0][6] ),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\partial_prod[2][2] ),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\partial_prod[0][0] ),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\partial_prod[1][2] ),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\partial_prod[0][13] ),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\partial_prod[0][2] ),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\partial_prod[2][1] ),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\partial_prod[1][10] ),
    .X(net116));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_56 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_215 ();
endmodule
